
module LASER_DW_mult_uns_3 ( a, b, product );
  input [6:0] a;
  input [6:0] b;
  output [13:0] product;
  wire   \a[0] , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111;
  assign product[0] = \a[0] ;
  assign \a[0]  = a[0];

  CLKXOR2X2 U54 ( .A(n84), .B(n86), .Y(product[4]) );
  XOR2X2 U55 ( .A(n103), .B(n102), .Y(n109) );
  CLKXOR2X2 U56 ( .A(n107), .B(n106), .Y(n108) );
  NOR2X2 U57 ( .A(n111), .B(n79), .Y(n107) );
  XOR2X4 U58 ( .A(n89), .B(n88), .Y(n91) );
  CLKXOR2X2 U59 ( .A(n93), .B(n94), .Y(n88) );
  AND2X2 U60 ( .A(n80), .B(\a[0] ), .Y(n83) );
  CLKINVX1 U61 ( .A(\a[0] ), .Y(n101) );
  BUFX8 U62 ( .A(a[3]), .Y(n80) );
  INVX3 U63 ( .A(a[1]), .Y(n111) );
  NAND2X1 U64 ( .A(n86), .B(n102), .Y(n92) );
  NOR2X1 U65 ( .A(n101), .B(n87), .Y(n94) );
  XOR2X1 U66 ( .A(n92), .B(n91), .Y(product[5]) );
  OR2X2 U67 ( .A(n96), .B(n101), .Y(n79) );
  XOR2X4 U68 ( .A(n100), .B(n99), .Y(product[6]) );
  NOR2BX2 U69 ( .AN(n90), .B(n96), .Y(n86) );
  INVX3 U70 ( .A(b[5]), .Y(n87) );
  XOR2X4 U71 ( .A(n109), .B(n108), .Y(product[3]) );
  OA21X2 U72 ( .A0(n92), .A1(n91), .B0(n90), .Y(n81) );
  INVX4 U73 ( .A(a[2]), .Y(n96) );
  NOR2XL U74 ( .A(n107), .B(n85), .Y(n84) );
  NOR2X2 U75 ( .A(n87), .B(n111), .Y(n93) );
  NOR2X4 U76 ( .A(n96), .B(n111), .Y(n82) );
  XOR2X1 U77 ( .A(n95), .B(n93), .Y(n89) );
  XNOR2X1 U78 ( .A(n81), .B(n93), .Y(n100) );
  NAND2X2 U79 ( .A(n83), .B(n82), .Y(n90) );
  XNOR2X4 U80 ( .A(n83), .B(n82), .Y(n85) );
  NAND2XL U81 ( .A(n95), .B(n94), .Y(n98) );
  CLKINVX1 U82 ( .A(n85), .Y(n102) );
  NAND2X1 U83 ( .A(a[1]), .B(n80), .Y(n95) );
  NAND2X1 U84 ( .A(n80), .B(n96), .Y(n97) );
  XOR2X1 U85 ( .A(n98), .B(n97), .Y(n99) );
  NOR2X1 U86 ( .A(n101), .B(n111), .Y(n110) );
  AO21X1 U87 ( .A0(\a[0] ), .A1(a[2]), .B0(n110), .Y(n103) );
  NAND2X1 U88 ( .A(a[2]), .B(a[1]), .Y(n105) );
  NAND2X1 U89 ( .A(\a[0] ), .B(n80), .Y(n104) );
  XOR2X1 U90 ( .A(n105), .B(n104), .Y(n106) );
  NOR2X1 U91 ( .A(n111), .B(n110), .Y(product[2]) );
endmodule


module LASER_DW_mult_uns_2 ( a, b, product );
  input [6:0] a;
  input [6:0] b;
  output [13:0] product;
  wire   \a[0] , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110;
  assign product[0] = \a[0] ;
  assign \a[0]  = a[0];

  INVX3 U54 ( .A(a[1]), .Y(n110) );
  AND2X2 U55 ( .A(a[3]), .B(\a[0] ), .Y(n81) );
  XOR2X2 U56 ( .A(n87), .B(n86), .Y(n89) );
  CLKBUFX3 U57 ( .A(n91), .Y(n79) );
  INVX3 U58 ( .A(n83), .Y(n101) );
  XOR2X1 U59 ( .A(n106), .B(n105), .Y(n107) );
  XOR2X2 U60 ( .A(n99), .B(n98), .Y(product[6]) );
  XOR2X1 U61 ( .A(n82), .B(n84), .Y(product[4]) );
  OAI21X2 U62 ( .A0(n90), .A1(n89), .B0(n88), .Y(n92) );
  INVX3 U63 ( .A(a[2]), .Y(n95) );
  NAND2X2 U64 ( .A(n84), .B(n101), .Y(n90) );
  NOR2BX2 U65 ( .AN(n88), .B(n95), .Y(n84) );
  XOR2X1 U66 ( .A(n90), .B(n89), .Y(product[5]) );
  NOR2XL U67 ( .A(n106), .B(n83), .Y(n82) );
  XNOR2X4 U68 ( .A(n81), .B(n80), .Y(n83) );
  XOR2X2 U69 ( .A(n108), .B(n107), .Y(product[3]) );
  XOR2X1 U70 ( .A(n92), .B(n79), .Y(n99) );
  NOR2X2 U71 ( .A(n95), .B(n110), .Y(n80) );
  CLKINVX1 U72 ( .A(\a[0] ), .Y(n100) );
  NOR3X1 U73 ( .A(n100), .B(n110), .C(n95), .Y(n106) );
  CLKINVX1 U74 ( .A(b[5]), .Y(n85) );
  NOR2X1 U75 ( .A(n100), .B(n85), .Y(n93) );
  NAND2X1 U76 ( .A(n81), .B(n80), .Y(n88) );
  NAND2X1 U77 ( .A(a[1]), .B(a[3]), .Y(n94) );
  NOR2X1 U78 ( .A(n85), .B(n110), .Y(n91) );
  XOR2X1 U79 ( .A(n94), .B(n79), .Y(n87) );
  XOR2X1 U80 ( .A(n79), .B(n93), .Y(n86) );
  NAND2X1 U81 ( .A(n94), .B(n93), .Y(n97) );
  NAND2X1 U82 ( .A(a[3]), .B(n95), .Y(n96) );
  XOR2X1 U83 ( .A(n97), .B(n96), .Y(n98) );
  NOR2X1 U84 ( .A(n100), .B(n110), .Y(n109) );
  AO21X1 U85 ( .A0(\a[0] ), .A1(a[2]), .B0(n109), .Y(n102) );
  XOR2X1 U86 ( .A(n102), .B(n101), .Y(n108) );
  NAND2X1 U87 ( .A(a[2]), .B(a[1]), .Y(n104) );
  NAND2X1 U88 ( .A(\a[0] ), .B(a[3]), .Y(n103) );
  XOR2X1 U89 ( .A(n104), .B(n103), .Y(n105) );
  NOR2X1 U90 ( .A(n110), .B(n109), .Y(product[2]) );
endmodule


module LASER_DW01_add_1 ( A, B, CI, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6;
  wire   [6:1] carry;

  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  AND2X2 U1 ( .A(B[2]), .B(A[2]), .Y(n1) );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[1]) );
  NAND2X2 U3 ( .A(B[4]), .B(carry[4]), .Y(n5) );
  NAND2X2 U4 ( .A(B[4]), .B(A[4]), .Y(n6) );
  XOR2XL U5 ( .A(A[4]), .B(B[4]), .Y(n3) );
  NAND2X2 U6 ( .A(A[4]), .B(carry[4]), .Y(n4) );
  XOR2X1 U7 ( .A(carry[4]), .B(n3), .Y(SUM[4]) );
  NAND3X2 U8 ( .A(n4), .B(n5), .C(n6), .Y(carry[5]) );
  XOR2XL U9 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  XOR2XL U10 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module LASER_DW_mult_uns_1 ( a, b, product );
  input [6:0] a;
  input [6:0] b;
  output [13:0] product;
  wire   \a[0] , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113;
  assign product[0] = \a[0] ;
  assign \a[0]  = a[0];

  CLKXOR2X4 U54 ( .A(n94), .B(n96), .Y(n89) );
  CLKXOR2X2 U55 ( .A(n109), .B(n108), .Y(n110) );
  XOR2X2 U56 ( .A(n85), .B(n87), .Y(product[4]) );
  NAND2X1 U57 ( .A(n87), .B(n104), .Y(n93) );
  NOR2BX2 U58 ( .AN(n91), .B(n98), .Y(n87) );
  XOR2X2 U59 ( .A(n105), .B(n104), .Y(n111) );
  INVX2 U60 ( .A(n86), .Y(n104) );
  INVX3 U61 ( .A(a[1]), .Y(n113) );
  CLKINVX1 U62 ( .A(\a[0] ), .Y(n103) );
  XOR2X2 U63 ( .A(n95), .B(n94), .Y(n102) );
  CLKINVX1 U64 ( .A(n83), .Y(n80) );
  AND2X2 U65 ( .A(a[3]), .B(\a[0] ), .Y(n84) );
  NAND2X1 U66 ( .A(n84), .B(n83), .Y(n91) );
  XOR2X2 U67 ( .A(n102), .B(n101), .Y(product[6]) );
  XOR2X4 U68 ( .A(n111), .B(n110), .Y(product[3]) );
  XOR2X4 U69 ( .A(n97), .B(n94), .Y(n90) );
  NOR2X2 U70 ( .A(n88), .B(n113), .Y(n94) );
  INVX8 U71 ( .A(a[2]), .Y(n98) );
  NOR2X1 U72 ( .A(n103), .B(n113), .Y(n112) );
  NAND2XL U73 ( .A(\a[0] ), .B(a[3]), .Y(n106) );
  NAND2XL U74 ( .A(a[3]), .B(n98), .Y(n99) );
  NAND2XL U75 ( .A(a[1]), .B(a[3]), .Y(n97) );
  INVX4 U76 ( .A(n84), .Y(n79) );
  NAND2X2 U77 ( .A(n84), .B(n83), .Y(n81) );
  NAND2X4 U78 ( .A(n79), .B(n80), .Y(n82) );
  NAND2X4 U79 ( .A(n81), .B(n82), .Y(n86) );
  NOR2XL U80 ( .A(n109), .B(n86), .Y(n85) );
  XOR2X1 U81 ( .A(n93), .B(n92), .Y(product[5]) );
  OAI21X1 U82 ( .A0(n93), .A1(n92), .B0(n91), .Y(n95) );
  NOR2X4 U83 ( .A(n98), .B(n113), .Y(n83) );
  NOR2XL U84 ( .A(n113), .B(n112), .Y(product[2]) );
  INVX3 U85 ( .A(b[5]), .Y(n88) );
  NOR2X1 U86 ( .A(n103), .B(n88), .Y(n96) );
  NOR3X1 U87 ( .A(n103), .B(n113), .C(n98), .Y(n109) );
  XOR2X1 U88 ( .A(n90), .B(n89), .Y(n92) );
  NAND2X1 U89 ( .A(n97), .B(n96), .Y(n100) );
  XOR2X1 U90 ( .A(n100), .B(n99), .Y(n101) );
  AO21X1 U91 ( .A0(\a[0] ), .A1(a[2]), .B0(n112), .Y(n105) );
  NAND2X1 U92 ( .A(a[2]), .B(a[1]), .Y(n107) );
  XOR2X1 U93 ( .A(n107), .B(n106), .Y(n108) );
endmodule


module LASER_DW_mult_uns_0 ( a, b, product );
  input [6:0] a;
  input [6:0] b;
  output [13:0] product;
  wire   \a[0] , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114;
  assign product[0] = \a[0] ;
  assign \a[0]  = a[0];

  NAND2XL U54 ( .A(n98), .B(n97), .Y(n101) );
  NOR2X2 U55 ( .A(n99), .B(n114), .Y(n85) );
  INVX3 U56 ( .A(a[1]), .Y(n114) );
  CLKINVX1 U57 ( .A(n95), .Y(n82) );
  NAND2X1 U58 ( .A(n86), .B(n85), .Y(n93) );
  AND2X2 U59 ( .A(a[3]), .B(\a[0] ), .Y(n86) );
  INVX3 U60 ( .A(a[2]), .Y(n99) );
  XOR2X1 U61 ( .A(n110), .B(n109), .Y(n111) );
  NOR2X2 U62 ( .A(n114), .B(n79), .Y(n110) );
  CLKINVX1 U63 ( .A(n80), .Y(n79) );
  NOR2BX1 U64 ( .AN(\a[0] ), .B(n99), .Y(n80) );
  NOR2BX1 U65 ( .AN(n93), .B(n99), .Y(n89) );
  XOR2X4 U66 ( .A(n112), .B(n111), .Y(product[3]) );
  NAND2X1 U67 ( .A(a[1]), .B(a[3]), .Y(n98) );
  NOR2X2 U68 ( .A(n90), .B(n114), .Y(n96) );
  INVX3 U69 ( .A(b[5]), .Y(n90) );
  XNOR2X2 U70 ( .A(n86), .B(n85), .Y(n88) );
  INVX1 U71 ( .A(\a[0] ), .Y(n104) );
  XOR2X4 U72 ( .A(n81), .B(n96), .Y(n103) );
  NAND2X2 U73 ( .A(n84), .B(n93), .Y(n81) );
  XOR2XL U74 ( .A(n95), .B(n94), .Y(product[5]) );
  NAND2X2 U75 ( .A(n89), .B(n105), .Y(n95) );
  XOR2X4 U76 ( .A(n103), .B(n102), .Y(product[6]) );
  NAND2X1 U77 ( .A(n82), .B(n83), .Y(n84) );
  XOR2X2 U78 ( .A(n92), .B(n91), .Y(n94) );
  CLKINVX1 U79 ( .A(n94), .Y(n83) );
  NOR2XL U80 ( .A(n110), .B(n88), .Y(n87) );
  INVX3 U81 ( .A(n88), .Y(n105) );
  NAND2XL U82 ( .A(\a[0] ), .B(a[3]), .Y(n107) );
  NOR2X1 U83 ( .A(n104), .B(n90), .Y(n97) );
  NAND2XL U84 ( .A(a[3]), .B(n99), .Y(n100) );
  AO21XL U85 ( .A0(\a[0] ), .A1(a[2]), .B0(n113), .Y(n106) );
  NAND2XL U86 ( .A(a[2]), .B(a[1]), .Y(n108) );
  XOR2X1 U87 ( .A(n87), .B(n89), .Y(product[4]) );
  XOR2X1 U88 ( .A(n98), .B(n96), .Y(n92) );
  XOR2X1 U89 ( .A(n96), .B(n97), .Y(n91) );
  XOR2X1 U90 ( .A(n101), .B(n100), .Y(n102) );
  NOR2X1 U91 ( .A(n104), .B(n114), .Y(n113) );
  XOR2X1 U92 ( .A(n106), .B(n105), .Y(n112) );
  XOR2X1 U93 ( .A(n108), .B(n107), .Y(n109) );
  NOR2X1 U94 ( .A(n114), .B(n113), .Y(product[2]) );
endmodule


module LASER_DW01_add_0 ( A, B, CI, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [6:1] carry;

  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  AND2X2 U1 ( .A(B[2]), .B(A[2]), .Y(n1) );
  AND2X2 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[1]) );
  XOR2XL U3 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module LASER ( CLK, RST, X, Y, C1X, C1Y, C2X, C2Y, DONE );
  input [3:0] X;
  input [3:0] Y;
  output [3:0] C1X;
  output [3:0] C1Y;
  output [3:0] C2X;
  output [3:0] C2Y;
  input CLK, RST;
  output DONE;
  wire   n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, \targetX[39][3] ,
         \targetX[39][2] , \targetX[39][1] , \targetX[39][0] ,
         \targetX[38][3] , \targetX[38][2] , \targetX[38][1] ,
         \targetX[38][0] , \targetX[37][3] , \targetX[37][2] ,
         \targetX[37][1] , \targetX[37][0] , \targetX[36][3] ,
         \targetX[36][2] , \targetX[36][1] , \targetX[36][0] ,
         \targetX[35][3] , \targetX[35][2] , \targetX[35][1] ,
         \targetX[35][0] , \targetX[34][3] , \targetX[34][2] ,
         \targetX[34][1] , \targetX[34][0] , \targetX[33][3] ,
         \targetX[33][2] , \targetX[33][1] , \targetX[33][0] ,
         \targetX[32][3] , \targetX[32][2] , \targetX[32][1] ,
         \targetX[32][0] , \targetX[15][3] , \targetX[15][0] ,
         \targetX[14][3] , \targetX[14][0] , \targetX[13][3] ,
         \targetX[13][0] , \targetX[12][3] , \targetX[12][0] ,
         \targetX[11][3] , \targetX[11][0] , \targetX[10][3] ,
         \targetX[10][0] , \targetX[9][3] , \targetX[9][0] , \targetX[8][3] ,
         \targetX[8][0] , \targetX[7][3] , \targetX[7][0] , \targetX[6][3] ,
         \targetX[6][0] , \targetX[5][3] , \targetX[5][0] , \targetX[4][3] ,
         \targetX[4][0] , \targetY[39][3] , \targetY[39][2] , \targetY[39][1] ,
         \targetY[39][0] , \targetY[38][3] , \targetY[38][2] ,
         \targetY[38][1] , \targetY[38][0] , \targetY[37][3] ,
         \targetY[37][2] , \targetY[37][1] , \targetY[37][0] ,
         \targetY[36][3] , \targetY[36][2] , \targetY[36][1] ,
         \targetY[36][0] , \targetY[35][3] , \targetY[35][2] ,
         \targetY[35][1] , \targetY[35][0] , \targetY[34][3] ,
         \targetY[34][2] , \targetY[34][1] , \targetY[34][0] ,
         \targetY[33][3] , \targetY[33][2] , \targetY[33][1] ,
         \targetY[33][0] , \targetY[32][3] , \targetY[32][2] ,
         \targetY[32][1] , \targetY[32][0] , \targetY[31][2] ,
         \targetY[31][0] , \targetY[30][2] , \targetY[30][0] ,
         \targetY[29][2] , \targetY[29][0] , \targetY[28][2] ,
         \targetY[28][0] , \targetY[27][2] , \targetY[27][1] ,
         \targetY[27][0] , \targetY[26][2] , \targetY[26][1] ,
         \targetY[26][0] , \targetY[25][2] , \targetY[25][1] ,
         \targetY[25][0] , \targetY[24][2] , \targetY[24][1] ,
         \targetY[24][0] , \targetY[23][0] , \targetY[22][0] ,
         \targetY[21][0] , \targetY[20][0] , \targetY[19][2] ,
         \targetY[19][1] , \targetY[19][0] , \targetY[18][2] ,
         \targetY[18][1] , \targetY[18][0] , \targetY[17][2] ,
         \targetY[17][1] , \targetY[17][0] , \targetY[16][2] ,
         \targetY[16][1] , \targetY[16][0] , \targetY[11][1] ,
         \targetY[10][1] , \targetY[9][1] , \targetY[8][1] , \targetY[7][1] ,
         \targetY[6][1] , \targetY[5][1] , \targetY[4][1] , \targetY[3][1] ,
         \targetY[2][1] , \targetY[1][1] , \targetY[0][1] , N826, N827, N828,
         N829, N830, N843, N844, N845, N846, N847, N903, N948, N949, N950,
         N951, N952, N965, N966, N967, N968, N969, N982, N983, N1020, N1021,
         N1022, N1023, optimise, N1049, N1050, N1051, N1052, N1053, N1130,
         N1131, N1132, N1133, N1134, n179, n185, n186, n187, n197, n198, n199,
         n200, n201, n202, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         N859, N858, N857, N856, N855, N853, N842, N841, N840, N839, N838,
         N836, N981, N980, N979, N978, N977, N975, N964, N963, N962, N961,
         N960, N958, \add_215/carry[5] , \add_215/carry[4] ,
         \add_215/carry[3] , \add_215/carry[2] , \r412/carry[5] ,
         \r412/carry[4] , \r412/carry[3] , \r412/carry[2] , \r406/carry[4] ,
         \r406/carry[3] , \r406/carry[2] , \r406/carry[1] , \r404/carry[4] ,
         \r404/carry[3] , \r404/carry[2] , \r404/carry[1] , \r401/carry[4] ,
         \r401/carry[3] , \r401/carry[2] , \r401/carry[1] , \r399/carry[4] ,
         \r399/carry[3] , \r399/carry[2] , \r399/carry[1] , n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568;
  wire   [5:0] count;
  wire   [6:0] len1;
  wire   [6:0] len2;
  wire   [2:0] state;
  wire   [2:0] nextState;
  wire   [5:0] covered;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31;

  LASER_DW_mult_uns_3 mult_36_2 ( .a({N847, N847, N847, N846, N845, N844, N843}), .b({N847, N847, N847, N846, N845, N844, N843}), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, N859, N858, N857, N856, N855, 
        SYNOPSYS_UNCONNECTED__7, N853}) );
  LASER_DW_mult_uns_2 mult_36 ( .a({N830, N830, N830, N829, N828, N827, N826}), 
        .b({N830, N830, N830, N829, N828, N827, N826}), .product({
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, N842, N841, N840, N839, N838, 
        SYNOPSYS_UNCONNECTED__15, N836}) );
  LASER_DW01_add_1 add_36 ( .A({N842, N841, N840, N839, N838, 1'b0, N836}), 
        .B({N859, N858, N857, N856, N855, 1'b0, N853}), .CI(1'b0), .SUM(len1)
         );
  LASER_DW_mult_uns_1 mult_37_2 ( .a({N969, N969, N969, N968, N967, N966, N965}), .b({N969, N969, N969, N968, N967, N966, N965}), .product({
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, N981, N980, N979, N978, N977, 
        SYNOPSYS_UNCONNECTED__23, N975}) );
  LASER_DW_mult_uns_0 mult_37 ( .a({N952, N952, N952, N951, N950, N949, N948}), 
        .b({N952, N952, N952, N951, N950, N949, N948}), .product({
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, N964, N963, N962, N961, N960, 
        SYNOPSYS_UNCONNECTED__31, N958}) );
  LASER_DW01_add_0 add_37 ( .A({N964, N963, N962, N961, N960, 1'b0, N958}), 
        .B({N981, N980, N979, N978, N977, 1'b0, N975}), .CI(1'b0), .SUM(len2)
         );
  DFFRX1 \yMax1_reg[1]  ( .D(n288), .CK(CLK), .RN(n1379), .QN(n1487) );
  DFFRX1 \yMax2_reg[1]  ( .D(n310), .CK(CLK), .RN(n1381), .QN(n1441) );
  DFFRX1 \covered_reg[3]  ( .D(n322), .CK(CLK), .RN(n1378), .Q(covered[3]), 
        .QN(n253) );
  DFFRX1 \covered_reg[4]  ( .D(n321), .CK(CLK), .RN(n1568), .Q(covered[4]), 
        .QN(n252) );
  DFFRX2 \covered_reg[5]  ( .D(n320), .CK(CLK), .RN(n1568), .Q(covered[5]), 
        .QN(n251) );
  EDFFX1 \targetX_reg[30][3]  ( .D(X[3]), .E(n223), .CK(CLK), .QN(n1132) );
  EDFFX1 \targetX_reg[30][2]  ( .D(X[2]), .E(n223), .CK(CLK), .QN(n1108) );
  EDFFX1 \targetY_reg[30][3]  ( .D(Y[3]), .E(n223), .CK(CLK), .QN(n1220) );
  EDFFX1 \targetX_reg[22][3]  ( .D(X[3]), .E(n222), .CK(CLK), .QN(n1156) );
  EDFFX1 \targetX_reg[22][2]  ( .D(X[2]), .E(n222), .CK(CLK), .QN(n1148) );
  EDFFX1 \targetY_reg[22][3]  ( .D(Y[3]), .E(n222), .CK(CLK), .QN(n1232) );
  EDFFX1 \targetX_reg[14][2]  ( .D(X[2]), .E(n221), .CK(CLK), .QN(n1196) );
  EDFFX1 \targetY_reg[14][3]  ( .D(Y[3]), .E(n221), .CK(CLK), .QN(n1208) );
  EDFFX1 \targetX_reg[6][2]  ( .D(X[2]), .E(n220), .CK(CLK), .QN(n1200) );
  EDFFX1 \targetY_reg[6][3]  ( .D(Y[3]), .E(n220), .CK(CLK), .QN(n1228) );
  EDFFX1 \targetY_reg[6][2]  ( .D(Y[2]), .E(n220), .CK(CLK), .QN(n1140) );
  EDFFX1 \targetX_reg[26][3]  ( .D(X[3]), .E(n213), .CK(CLK), .QN(n1248) );
  EDFFX1 \targetX_reg[26][2]  ( .D(X[2]), .E(n213), .CK(CLK), .QN(n1168) );
  EDFFX1 \targetY_reg[26][3]  ( .D(Y[3]), .E(n213), .CK(CLK), .QN(n1216) );
  EDFFX1 \targetX_reg[18][3]  ( .D(X[3]), .E(n212), .CK(CLK), .QN(n1240) );
  EDFFX1 \targetX_reg[18][2]  ( .D(X[2]), .E(n212), .CK(CLK), .QN(n1128) );
  EDFFX1 \targetY_reg[18][3]  ( .D(Y[3]), .E(n212), .CK(CLK), .QN(n1212) );
  EDFFX1 \targetX_reg[10][2]  ( .D(X[2]), .E(n211), .CK(CLK), .QN(n1204) );
  EDFFX1 \targetY_reg[10][3]  ( .D(Y[3]), .E(n211), .CK(CLK), .QN(n1244) );
  EDFFX1 \targetX_reg[2][3]  ( .D(X[3]), .E(n210), .CK(CLK), .QN(n1236) );
  EDFFX1 \targetX_reg[2][2]  ( .D(X[2]), .E(n210), .CK(CLK), .QN(n1152) );
  EDFFX1 \targetX_reg[2][1]  ( .D(X[1]), .E(n210), .CK(CLK), .QN(n1116) );
  EDFFX1 \targetY_reg[2][3]  ( .D(Y[3]), .E(n210), .CK(CLK), .QN(n1224) );
  EDFFX1 \targetY_reg[2][2]  ( .D(Y[2]), .E(n210), .CK(CLK), .QN(n1124) );
  EDFFX1 \targetX_reg[31][3]  ( .D(X[3]), .E(n243), .CK(CLK), .QN(n1134) );
  EDFFX1 \targetX_reg[31][2]  ( .D(X[2]), .E(n243), .CK(CLK), .QN(n1110) );
  EDFFX1 \targetY_reg[31][3]  ( .D(Y[3]), .E(n243), .CK(CLK), .QN(n1222) );
  EDFFX1 \targetX_reg[23][3]  ( .D(X[3]), .E(n242), .CK(CLK), .QN(n1158) );
  EDFFX1 \targetX_reg[23][2]  ( .D(X[2]), .E(n242), .CK(CLK), .QN(n1150) );
  EDFFX1 \targetY_reg[23][3]  ( .D(Y[3]), .E(n242), .CK(CLK), .QN(n1234) );
  EDFFX1 \targetX_reg[15][2]  ( .D(X[2]), .E(n241), .CK(CLK), .QN(n1198) );
  EDFFX1 \targetY_reg[15][3]  ( .D(Y[3]), .E(n241), .CK(CLK), .QN(n1210) );
  EDFFX1 \targetY_reg[15][2]  ( .D(Y[2]), .E(n241), .CK(CLK), .QN(n1106) );
  EDFFX1 \targetX_reg[7][2]  ( .D(X[2]), .E(n240), .CK(CLK), .QN(n1202) );
  EDFFX1 \targetY_reg[7][3]  ( .D(Y[3]), .E(n240), .CK(CLK), .QN(n1230) );
  EDFFX1 \targetX_reg[27][3]  ( .D(X[3]), .E(n238), .CK(CLK), .QN(n1250) );
  EDFFX1 \targetX_reg[27][2]  ( .D(X[2]), .E(n238), .CK(CLK), .QN(n1170) );
  EDFFX1 \targetY_reg[27][3]  ( .D(Y[3]), .E(n238), .CK(CLK), .QN(n1218) );
  EDFFX1 \targetX_reg[19][3]  ( .D(X[3]), .E(n237), .CK(CLK), .QN(n1242) );
  EDFFX1 \targetX_reg[19][2]  ( .D(X[2]), .E(n237), .CK(CLK), .QN(n1130) );
  EDFFX1 \targetY_reg[19][3]  ( .D(Y[3]), .E(n237), .CK(CLK), .QN(n1214) );
  EDFFX1 \targetX_reg[11][2]  ( .D(X[2]), .E(n236), .CK(CLK), .QN(n1206) );
  EDFFX1 \targetX_reg[11][1]  ( .D(X[1]), .E(n236), .CK(CLK), .QN(n1194) );
  EDFFX1 \targetY_reg[11][3]  ( .D(Y[3]), .E(n236), .CK(CLK), .QN(n1246) );
  EDFFX1 \targetY_reg[11][2]  ( .D(Y[2]), .E(n236), .CK(CLK), .QN(n1166) );
  EDFFX1 \targetX_reg[3][3]  ( .D(X[3]), .E(n235), .CK(CLK), .QN(n1238) );
  EDFFX1 \targetX_reg[3][2]  ( .D(X[2]), .E(n235), .CK(CLK), .QN(n1154) );
  EDFFX1 \targetY_reg[3][3]  ( .D(Y[3]), .E(n235), .CK(CLK), .QN(n1226) );
  EDFFX1 \targetX_reg[28][3]  ( .D(X[3]), .E(n218), .CK(CLK), .QN(n1131) );
  EDFFX1 \targetX_reg[28][2]  ( .D(X[2]), .E(n218), .CK(CLK), .QN(n1107) );
  EDFFX1 \targetY_reg[28][3]  ( .D(Y[3]), .E(n218), .CK(CLK), .QN(n1219) );
  EDFFX1 \targetX_reg[20][3]  ( .D(X[3]), .E(n217), .CK(CLK), .QN(n1155) );
  EDFFX1 \targetX_reg[20][2]  ( .D(X[2]), .E(n217), .CK(CLK), .QN(n1147) );
  EDFFX1 \targetY_reg[20][3]  ( .D(Y[3]), .E(n217), .CK(CLK), .QN(n1231) );
  EDFFX1 \targetX_reg[12][2]  ( .D(X[2]), .E(n216), .CK(CLK), .QN(n1195) );
  EDFFX1 \targetY_reg[12][3]  ( .D(Y[3]), .E(n216), .CK(CLK), .QN(n1207) );
  EDFFX1 \targetX_reg[4][2]  ( .D(X[2]), .E(n215), .CK(CLK), .QN(n1199) );
  EDFFX1 \targetY_reg[4][3]  ( .D(Y[3]), .E(n215), .CK(CLK), .QN(n1227) );
  EDFFX1 \targetX_reg[24][3]  ( .D(X[3]), .E(n208), .CK(CLK), .QN(n1247) );
  EDFFX1 \targetX_reg[24][2]  ( .D(X[2]), .E(n208), .CK(CLK), .QN(n1167) );
  EDFFX1 \targetX_reg[24][1]  ( .D(X[1]), .E(n208), .CK(CLK), .QN(n1159) );
  EDFFX1 \targetX_reg[24][0]  ( .D(X[0]), .E(n208), .CK(CLK), .QN(n1078) );
  EDFFX1 \targetY_reg[24][3]  ( .D(Y[3]), .E(n208), .CK(CLK), .QN(n1215) );
  EDFFX1 \targetX_reg[16][3]  ( .D(X[3]), .E(n207), .CK(CLK), .QN(n1239) );
  EDFFX1 \targetX_reg[16][2]  ( .D(X[2]), .E(n207), .CK(CLK), .QN(n1127) );
  EDFFX1 \targetY_reg[16][3]  ( .D(Y[3]), .E(n207), .CK(CLK), .QN(n1211) );
  EDFFX1 \targetX_reg[8][2]  ( .D(X[2]), .E(n206), .CK(CLK), .QN(n1203) );
  EDFFX1 \targetY_reg[8][3]  ( .D(Y[3]), .E(n206), .CK(CLK), .QN(n1243) );
  EDFFX1 \targetX_reg[0][3]  ( .D(X[3]), .E(n205), .CK(CLK), .QN(n1235) );
  EDFFX1 \targetX_reg[0][2]  ( .D(X[2]), .E(n205), .CK(CLK), .QN(n1151) );
  EDFFX1 \targetY_reg[0][3]  ( .D(Y[3]), .E(n205), .CK(CLK), .QN(n1223) );
  EDFFX1 \targetX_reg[29][3]  ( .D(X[3]), .E(n233), .CK(CLK), .QN(n1133) );
  EDFFX1 \targetX_reg[29][2]  ( .D(X[2]), .E(n233), .CK(CLK), .QN(n1109) );
  EDFFX1 \targetY_reg[29][3]  ( .D(Y[3]), .E(n233), .CK(CLK), .QN(n1221) );
  EDFFX1 \targetX_reg[21][3]  ( .D(X[3]), .E(n232), .CK(CLK), .QN(n1157) );
  EDFFX1 \targetX_reg[21][2]  ( .D(X[2]), .E(n232), .CK(CLK), .QN(n1149) );
  EDFFX1 \targetY_reg[21][3]  ( .D(Y[3]), .E(n232), .CK(CLK), .QN(n1233) );
  EDFFX1 \targetY_reg[21][2]  ( .D(Y[2]), .E(n232), .CK(CLK), .QN(n1145) );
  EDFFX1 \targetX_reg[13][2]  ( .D(X[2]), .E(n231), .CK(CLK), .QN(n1197) );
  EDFFX1 \targetY_reg[13][3]  ( .D(Y[3]), .E(n231), .CK(CLK), .QN(n1209) );
  EDFFX1 \targetX_reg[5][2]  ( .D(X[2]), .E(n230), .CK(CLK), .QN(n1201) );
  EDFFX1 \targetY_reg[5][3]  ( .D(Y[3]), .E(n230), .CK(CLK), .QN(n1229) );
  EDFFX1 \targetX_reg[25][3]  ( .D(X[3]), .E(n228), .CK(CLK), .QN(n1249) );
  EDFFX1 \targetX_reg[25][2]  ( .D(X[2]), .E(n228), .CK(CLK), .QN(n1169) );
  EDFFX1 \targetY_reg[25][3]  ( .D(Y[3]), .E(n228), .CK(CLK), .QN(n1217) );
  EDFFX1 \targetX_reg[17][3]  ( .D(X[3]), .E(n227), .CK(CLK), .QN(n1241) );
  EDFFX1 \targetX_reg[17][2]  ( .D(X[2]), .E(n227), .CK(CLK), .QN(n1129) );
  EDFFX1 \targetX_reg[17][1]  ( .D(X[1]), .E(n227), .CK(CLK), .QN(n1121) );
  EDFFX1 \targetX_reg[17][0]  ( .D(X[0]), .E(n227), .CK(CLK), .QN(n1072) );
  EDFFX1 \targetY_reg[17][3]  ( .D(Y[3]), .E(n227), .CK(CLK), .QN(n1213) );
  EDFFX1 \targetX_reg[9][1]  ( .D(X[1]), .E(n226), .CK(CLK), .QN(n1193) );
  EDFFX1 \targetY_reg[9][3]  ( .D(Y[3]), .E(n226), .CK(CLK), .QN(n1245) );
  EDFFX1 \targetX_reg[1][3]  ( .D(X[3]), .E(n225), .CK(CLK), .QN(n1237) );
  EDFFX1 \targetX_reg[1][2]  ( .D(X[2]), .E(n225), .CK(CLK), .QN(n1153) );
  EDFFX1 \targetY_reg[1][3]  ( .D(Y[3]), .E(n225), .CK(CLK), .QN(n1225) );
  DFFRX1 \covered_reg[0]  ( .D(n325), .CK(CLK), .RN(n1378), .Q(covered[0]), 
        .QN(n256) );
  DFFRX1 \covered_reg[1]  ( .D(n324), .CK(CLK), .RN(n1378), .Q(covered[1]), 
        .QN(n255) );
  DFFRX1 \covered_reg[2]  ( .D(n323), .CK(CLK), .RN(n1378), .Q(covered[2]), 
        .QN(n254) );
  DFFRX1 \state_reg[0]  ( .D(nextState[0]), .CK(CLK), .RN(n1378), .Q(state[0]), 
        .QN(n1044) );
  DFFRX2 \state_reg[1]  ( .D(nextState[1]), .CK(CLK), .RN(n1378), .Q(state[1]), 
        .QN(n1046) );
  EDFFX1 \targetX_reg[2][0]  ( .D(X[0]), .E(n210), .CK(CLK), .QN(n1112) );
  EDFFX1 \targetY_reg[2][0]  ( .D(Y[0]), .E(n210), .CK(CLK), .QN(n1087) );
  EDFFX1 \targetY_reg[11][0]  ( .D(Y[0]), .E(n236), .CK(CLK), .QN(n1097) );
  ADDHXL \add_215/U1_1_4  ( .A(covered[4]), .B(\add_215/carry[4] ), .CO(
        \add_215/carry[5] ), .S(N1133) );
  ADDHXL \r412/U1_1_4  ( .A(count[4]), .B(\r412/carry[4] ), .CO(
        \r412/carry[5] ), .S(N1052) );
  ADDHXL \add_215/U1_1_3  ( .A(covered[3]), .B(\add_215/carry[3] ), .CO(
        \add_215/carry[4] ), .S(N1132) );
  ADDHXL \add_215/U1_1_2  ( .A(covered[2]), .B(\add_215/carry[2] ), .CO(
        \add_215/carry[3] ), .S(N1131) );
  ADDHXL \add_215/U1_1_1  ( .A(covered[1]), .B(covered[0]), .CO(
        \add_215/carry[2] ), .S(N1130) );
  ADDHXL \r412/U1_1_3  ( .A(count[3]), .B(\r412/carry[3] ), .CO(
        \r412/carry[4] ), .S(N1051) );
  TLATX1 \nextState_reg[0]  ( .G(N1020), .D(N1021), .Q(nextState[0]) );
  TLATX1 \nextState_reg[2]  ( .G(N1020), .D(N1023), .Q(nextState[2]) );
  TLATX1 \nextState_reg[1]  ( .G(N1020), .D(N1022), .Q(nextState[1]) );
  ADDHXL \r412/U1_1_1  ( .A(n1039), .B(n1374), .CO(\r412/carry[2] ), .S(N1049)
         );
  ADDHXL \r412/U1_1_2  ( .A(count[2]), .B(\r412/carry[2] ), .CO(
        \r412/carry[3] ), .S(N1050) );
  DFFRX4 \count_reg[0]  ( .D(n331), .CK(CLK), .RN(n1568), .Q(count[0]), .QN(
        n262) );
  DFFRHQX4 \count_reg[1]  ( .D(n330), .CK(CLK), .RN(n1379), .Q(n1061) );
  DFFRX1 \C1X_reg[0]  ( .D(n296), .CK(CLK), .RN(n1380), .Q(n1574), .QN(n269)
         );
  DFFRX1 \C2X_reg[0]  ( .D(n334), .CK(CLK), .RN(n1378), .Q(n1582), .QN(n276)
         );
  DFFRX1 \C2Y_reg[0]  ( .D(n313), .CK(CLK), .RN(n1381), .Q(n1586), .QN(n250)
         );
  DFFRX1 \C1X_reg[1]  ( .D(n294), .CK(CLK), .RN(n1380), .Q(n1573), .QN(n268)
         );
  DFFRX1 \C2X_reg[1]  ( .D(n316), .CK(CLK), .RN(n1380), .Q(n1581), .QN(n275)
         );
  DFFRX1 \C1Y_reg[2]  ( .D(n287), .CK(CLK), .RN(n1379), .Q(n1576), .QN(n271)
         );
  DFFRX1 \C2Y_reg[1]  ( .D(n311), .CK(CLK), .RN(n1381), .Q(n1585), .QN(n249)
         );
  DFFRX1 \C1X_reg[2]  ( .D(n292), .CK(CLK), .RN(n1380), .Q(n1572), .QN(n267)
         );
  DFFRX1 \C1X_reg[3]  ( .D(n298), .CK(CLK), .RN(n1380), .Q(n1571), .QN(n266)
         );
  DFFRX1 \C1Y_reg[3]  ( .D(n299), .CK(CLK), .RN(n1379), .Q(n1575), .QN(n270)
         );
  DFFRX1 \C2Y_reg[2]  ( .D(n309), .CK(CLK), .RN(n1381), .Q(n1584), .QN(n248)
         );
  DFFRX1 \C2Y_reg[3]  ( .D(n317), .CK(CLK), .RN(n1381), .Q(n1583), .QN(n247)
         );
  DFFRX1 \C2X_reg[3]  ( .D(n333), .CK(CLK), .RN(n1381), .Q(n1579), .QN(n204)
         );
  DFFRX1 \C1Y_reg[1]  ( .D(n289), .CK(CLK), .RN(n1379), .Q(n1577), .QN(n272)
         );
  DFFRX1 \C1Y_reg[0]  ( .D(n291), .CK(CLK), .RN(n1379), .Q(n1578), .QN(n273)
         );
  DFFRX1 \C2X_reg[2]  ( .D(n314), .CK(CLK), .RN(n1381), .Q(n1580), .QN(n274)
         );
  DFFRX1 DONE_reg ( .D(n332), .CK(CLK), .RN(n1379), .Q(n1587), .QN(n179) );
  ADDFHX2 \r406/U2_2  ( .A(C2Y[2]), .B(n1042), .CI(\r406/carry[2] ), .CO(
        \r406/carry[3] ), .S(N967) );
  ADDFHX2 \r406/U2_1  ( .A(C2Y[1]), .B(n1389), .CI(\r406/carry[1] ), .CO(
        \r406/carry[2] ), .S(N966) );
  ADDFHX2 \r399/U2_1  ( .A(C1X[1]), .B(n1384), .CI(\r399/carry[1] ), .CO(
        \r399/carry[2] ), .S(N827) );
  ADDFHX4 \r406/U2_3  ( .A(n1583), .B(n1040), .CI(\r406/carry[3] ), .CO(
        \r406/carry[4] ), .S(N968) );
  ADDFHX2 \r401/U2_2  ( .A(n1576), .B(n1042), .CI(\r401/carry[2] ), .CO(
        \r401/carry[3] ), .S(N845) );
  ADDFHX4 \r404/U2_1  ( .A(n1581), .B(n1388), .CI(\r404/carry[1] ), .CO(
        \r404/carry[2] ), .S(N949) );
  ADDFHX4 \r404/U2_3  ( .A(n1579), .B(n1385), .CI(\r404/carry[3] ), .CO(
        \r404/carry[4] ), .S(N951) );
  ADDFHX2 \r401/U2_1  ( .A(n1577), .B(n1389), .CI(\r401/carry[1] ), .CO(
        \r401/carry[2] ), .S(N844) );
  DFFSX1 doingC1_reg ( .D(n301), .CK(CLK), .SN(n1568), .Q(n1567), .QN(n1455)
         );
  EDFFXL \targetY_reg[33][1]  ( .D(Y[1]), .E(n229), .CK(CLK), .Q(
        \targetY[33][1] ) );
  EDFFXL \targetY_reg[33][0]  ( .D(Y[0]), .E(n229), .CK(CLK), .Q(
        \targetY[33][0] ) );
  EDFFXL \targetX_reg[33][1]  ( .D(X[1]), .E(n229), .CK(CLK), .Q(
        \targetX[33][1] ) );
  EDFFXL \targetX_reg[33][0]  ( .D(X[0]), .E(n229), .CK(CLK), .Q(
        \targetX[33][0] ) );
  EDFFXL \targetY_reg[37][2]  ( .D(Y[2]), .E(n234), .CK(CLK), .Q(
        \targetY[37][2] ) );
  EDFFXL \targetY_reg[37][1]  ( .D(Y[1]), .E(n234), .CK(CLK), .Q(
        \targetY[37][1] ) );
  EDFFXL \targetY_reg[37][0]  ( .D(Y[0]), .E(n234), .CK(CLK), .Q(
        \targetY[37][0] ) );
  EDFFXL \targetX_reg[37][1]  ( .D(X[1]), .E(n234), .CK(CLK), .Q(
        \targetX[37][1] ) );
  EDFFXL \targetX_reg[37][0]  ( .D(X[0]), .E(n234), .CK(CLK), .Q(
        \targetX[37][0] ) );
  EDFFXL \targetY_reg[38][2]  ( .D(Y[2]), .E(n224), .CK(CLK), .Q(
        \targetY[38][2] ) );
  EDFFXL \targetY_reg[38][1]  ( .D(Y[1]), .E(n224), .CK(CLK), .Q(
        \targetY[38][1] ) );
  EDFFXL \targetY_reg[38][0]  ( .D(Y[0]), .E(n224), .CK(CLK), .Q(
        \targetY[38][0] ) );
  EDFFXL \targetY_reg[36][2]  ( .D(Y[2]), .E(n219), .CK(CLK), .Q(
        \targetY[36][2] ) );
  EDFFXL \targetY_reg[36][1]  ( .D(Y[1]), .E(n219), .CK(CLK), .Q(
        \targetY[36][1] ) );
  EDFFXL \targetY_reg[36][0]  ( .D(Y[0]), .E(n219), .CK(CLK), .Q(
        \targetY[36][0] ) );
  EDFFXL \targetX_reg[38][1]  ( .D(X[1]), .E(n224), .CK(CLK), .Q(
        \targetX[38][1] ) );
  EDFFXL \targetX_reg[38][0]  ( .D(X[0]), .E(n224), .CK(CLK), .Q(
        \targetX[38][0] ) );
  EDFFXL \targetX_reg[36][1]  ( .D(X[1]), .E(n219), .CK(CLK), .Q(
        \targetX[36][1] ) );
  EDFFXL \targetX_reg[36][0]  ( .D(X[0]), .E(n219), .CK(CLK), .Q(
        \targetX[36][0] ) );
  EDFFXL \targetY_reg[34][2]  ( .D(Y[2]), .E(n214), .CK(CLK), .Q(
        \targetY[34][2] ) );
  EDFFXL \targetY_reg[34][1]  ( .D(Y[1]), .E(n214), .CK(CLK), .Q(
        \targetY[34][1] ) );
  EDFFXL \targetY_reg[34][0]  ( .D(Y[0]), .E(n214), .CK(CLK), .Q(
        \targetY[34][0] ) );
  EDFFXL \targetY_reg[32][2]  ( .D(Y[2]), .E(n209), .CK(CLK), .Q(
        \targetY[32][2] ) );
  EDFFXL \targetY_reg[32][1]  ( .D(Y[1]), .E(n209), .CK(CLK), .Q(
        \targetY[32][1] ) );
  EDFFXL \targetY_reg[32][0]  ( .D(Y[0]), .E(n209), .CK(CLK), .Q(
        \targetY[32][0] ) );
  EDFFXL \targetX_reg[34][2]  ( .D(X[2]), .E(n214), .CK(CLK), .Q(
        \targetX[34][2] ) );
  EDFFXL \targetX_reg[34][1]  ( .D(X[1]), .E(n214), .CK(CLK), .Q(
        \targetX[34][1] ) );
  EDFFXL \targetX_reg[32][1]  ( .D(X[1]), .E(n209), .CK(CLK), .Q(
        \targetX[32][1] ) );
  EDFFXL \targetX_reg[32][0]  ( .D(X[0]), .E(n209), .CK(CLK), .Q(
        \targetX[32][0] ) );
  EDFFXL \targetY_reg[33][2]  ( .D(Y[2]), .E(n229), .CK(CLK), .Q(
        \targetY[33][2] ) );
  EDFFXL \targetY_reg[31][2]  ( .D(Y[2]), .E(n243), .CK(CLK), .Q(
        \targetY[31][2] ) );
  EDFFXL \targetY_reg[31][0]  ( .D(Y[0]), .E(n243), .CK(CLK), .Q(
        \targetY[31][0] ) );
  EDFFXL \targetY_reg[23][0]  ( .D(Y[0]), .E(n242), .CK(CLK), .Q(
        \targetY[23][0] ) );
  EDFFXL \targetY_reg[7][1]  ( .D(Y[1]), .E(n240), .CK(CLK), .Q(
        \targetY[7][1] ) );
  EDFFXL \targetX_reg[7][0]  ( .D(X[0]), .E(n240), .CK(CLK), .Q(
        \targetX[7][0] ) );
  EDFFXL \targetY_reg[29][2]  ( .D(Y[2]), .E(n233), .CK(CLK), .Q(
        \targetY[29][2] ) );
  EDFFXL \targetY_reg[29][0]  ( .D(Y[0]), .E(n233), .CK(CLK), .Q(
        \targetY[29][0] ) );
  EDFFXL \targetY_reg[25][2]  ( .D(Y[2]), .E(n228), .CK(CLK), .Q(
        \targetY[25][2] ) );
  EDFFXL \targetY_reg[25][1]  ( .D(Y[1]), .E(n228), .CK(CLK), .Q(
        \targetY[25][1] ) );
  EDFFXL \targetY_reg[25][0]  ( .D(Y[0]), .E(n228), .CK(CLK), .Q(
        \targetY[25][0] ) );
  EDFFXL \targetY_reg[9][1]  ( .D(Y[1]), .E(n226), .CK(CLK), .Q(
        \targetY[9][1] ) );
  EDFFXL \targetY_reg[5][1]  ( .D(Y[1]), .E(n230), .CK(CLK), .Q(
        \targetY[5][1] ) );
  EDFFXL \targetY_reg[1][1]  ( .D(Y[1]), .E(n225), .CK(CLK), .Q(
        \targetY[1][1] ) );
  EDFFXL \targetX_reg[13][0]  ( .D(X[0]), .E(n231), .CK(CLK), .Q(
        \targetX[13][0] ) );
  EDFFXL \targetX_reg[9][0]  ( .D(X[0]), .E(n226), .CK(CLK), .Q(
        \targetX[9][0] ) );
  EDFFXL \targetX_reg[5][0]  ( .D(X[0]), .E(n230), .CK(CLK), .Q(
        \targetX[5][0] ) );
  EDFFXL \targetY_reg[30][2]  ( .D(Y[2]), .E(n223), .CK(CLK), .Q(
        \targetY[30][2] ) );
  EDFFXL \targetY_reg[30][0]  ( .D(Y[0]), .E(n223), .CK(CLK), .Q(
        \targetY[30][0] ) );
  EDFFXL \targetY_reg[22][0]  ( .D(Y[0]), .E(n222), .CK(CLK), .Q(
        \targetY[22][0] ) );
  EDFFXL \targetY_reg[20][0]  ( .D(Y[0]), .E(n217), .CK(CLK), .Q(
        \targetY[20][0] ) );
  EDFFXL \targetY_reg[4][1]  ( .D(Y[1]), .E(n215), .CK(CLK), .Q(
        \targetY[4][1] ) );
  EDFFXL \targetX_reg[14][0]  ( .D(X[0]), .E(n221), .CK(CLK), .Q(
        \targetX[14][0] ) );
  EDFFXL \targetX_reg[12][0]  ( .D(X[0]), .E(n216), .CK(CLK), .Q(
        \targetX[12][0] ) );
  EDFFXL \targetX_reg[4][0]  ( .D(X[0]), .E(n215), .CK(CLK), .Q(
        \targetX[4][0] ) );
  EDFFXL \targetY_reg[27][2]  ( .D(Y[2]), .E(n238), .CK(CLK), .Q(
        \targetY[27][2] ) );
  EDFFXL \targetY_reg[27][1]  ( .D(Y[1]), .E(n238), .CK(CLK), .Q(
        \targetY[27][1] ) );
  EDFFXL \targetY_reg[27][0]  ( .D(Y[0]), .E(n238), .CK(CLK), .Q(
        \targetY[27][0] ) );
  EDFFXL \targetY_reg[19][2]  ( .D(Y[2]), .E(n237), .CK(CLK), .Q(
        \targetY[19][2] ) );
  EDFFXL \targetY_reg[19][1]  ( .D(Y[1]), .E(n237), .CK(CLK), .Q(
        \targetY[19][1] ) );
  EDFFXL \targetY_reg[19][0]  ( .D(Y[0]), .E(n237), .CK(CLK), .Q(
        \targetY[19][0] ) );
  EDFFXL \targetY_reg[3][1]  ( .D(Y[1]), .E(n235), .CK(CLK), .Q(
        \targetY[3][1] ) );
  EDFFXL \targetY_reg[26][2]  ( .D(Y[2]), .E(n213), .CK(CLK), .Q(
        \targetY[26][2] ) );
  EDFFXL \targetY_reg[26][1]  ( .D(Y[1]), .E(n213), .CK(CLK), .Q(
        \targetY[26][1] ) );
  EDFFXL \targetY_reg[26][0]  ( .D(Y[0]), .E(n213), .CK(CLK), .Q(
        \targetY[26][0] ) );
  EDFFXL \targetY_reg[18][2]  ( .D(Y[2]), .E(n212), .CK(CLK), .Q(
        \targetY[18][2] ) );
  EDFFXL \targetY_reg[18][1]  ( .D(Y[1]), .E(n212), .CK(CLK), .Q(
        \targetY[18][1] ) );
  EDFFXL \targetY_reg[18][0]  ( .D(Y[0]), .E(n212), .CK(CLK), .Q(
        \targetY[18][0] ) );
  EDFFXL \targetY_reg[16][2]  ( .D(Y[2]), .E(n207), .CK(CLK), .Q(
        \targetY[16][2] ) );
  EDFFXL \targetY_reg[16][1]  ( .D(Y[1]), .E(n207), .CK(CLK), .Q(
        \targetY[16][1] ) );
  EDFFXL \targetY_reg[16][0]  ( .D(Y[0]), .E(n207), .CK(CLK), .Q(
        \targetY[16][0] ) );
  EDFFXL \targetY_reg[10][1]  ( .D(Y[1]), .E(n211), .CK(CLK), .Q(
        \targetY[10][1] ) );
  EDFFXL \targetY_reg[8][1]  ( .D(Y[1]), .E(n206), .CK(CLK), .Q(
        \targetY[8][1] ) );
  EDFFXL \targetY_reg[0][1]  ( .D(Y[1]), .E(n205), .CK(CLK), .Q(
        \targetY[0][1] ) );
  EDFFXL \targetX_reg[10][0]  ( .D(X[0]), .E(n211), .CK(CLK), .Q(
        \targetX[10][0] ) );
  EDFFXL \targetX_reg[8][0]  ( .D(X[0]), .E(n206), .CK(CLK), .Q(
        \targetX[8][0] ) );
  EDFFXL \targetX_reg[15][0]  ( .D(X[0]), .E(n241), .CK(CLK), .Q(
        \targetX[15][0] ) );
  EDFFXL \targetX_reg[6][0]  ( .D(X[0]), .E(n220), .CK(CLK), .Q(
        \targetX[6][0] ) );
  EDFFXL \targetY_reg[15][0]  ( .D(Y[0]), .E(n241), .CK(CLK), .QN(n1093) );
  EDFFXL \targetX_reg[15][1]  ( .D(X[1]), .E(n241), .CK(CLK), .QN(n1186) );
  EDFFXL \targetY_reg[31][1]  ( .D(Y[1]), .E(n243), .CK(CLK), .QN(n1182) );
  EDFFXL \targetY_reg[23][2]  ( .D(Y[2]), .E(n242), .CK(CLK), .QN(n1146) );
  EDFFXL \targetY_reg[23][1]  ( .D(Y[1]), .E(n242), .CK(CLK), .QN(n1178) );
  EDFFXL \targetY_reg[7][2]  ( .D(Y[2]), .E(n240), .CK(CLK), .QN(n1142) );
  EDFFXL \targetY_reg[7][0]  ( .D(Y[0]), .E(n240), .CK(CLK), .QN(n1085) );
  EDFFXL \targetX_reg[31][1]  ( .D(X[1]), .E(n243), .CK(CLK), .QN(n1102) );
  EDFFXL \targetX_reg[31][0]  ( .D(X[0]), .E(n243), .CK(CLK), .QN(n1077) );
  EDFFXL \targetX_reg[23][1]  ( .D(X[1]), .E(n242), .CK(CLK), .QN(n1138) );
  EDFFXL \targetX_reg[23][0]  ( .D(X[0]), .E(n242), .CK(CLK), .QN(n1069) );
  EDFFXL \targetX_reg[7][1]  ( .D(X[1]), .E(n240), .CK(CLK), .QN(n1190) );
  EDFFXL \targetY_reg[21][1]  ( .D(Y[1]), .E(n232), .CK(CLK), .QN(n1177) );
  EDFFXL \targetX_reg[21][1]  ( .D(X[1]), .E(n232), .CK(CLK), .QN(n1137) );
  EDFFXL \targetY_reg[28][1]  ( .D(Y[1]), .E(n218), .CK(CLK), .QN(n1179) );
  EDFFXL \targetY_reg[6][0]  ( .D(Y[0]), .E(n220), .CK(CLK), .QN(n1083) );
  EDFFXL \targetX_reg[28][1]  ( .D(X[1]), .E(n218), .CK(CLK), .QN(n1099) );
  EDFFXL \targetX_reg[6][1]  ( .D(X[1]), .E(n220), .CK(CLK), .QN(n1188) );
  EDFFXL \targetY_reg[29][1]  ( .D(Y[1]), .E(n233), .CK(CLK), .QN(n1181) );
  EDFFXL \targetY_reg[13][2]  ( .D(Y[2]), .E(n231), .CK(CLK), .QN(n1105) );
  EDFFXL \targetY_reg[13][1]  ( .D(Y[1]), .E(n231), .CK(CLK), .QN(n1173) );
  EDFFXL \targetY_reg[13][0]  ( .D(Y[0]), .E(n231), .CK(CLK), .QN(n1092) );
  EDFFXL \targetY_reg[9][2]  ( .D(Y[2]), .E(n226), .CK(CLK), .QN(n1165) );
  EDFFXL \targetY_reg[9][0]  ( .D(Y[0]), .E(n226), .CK(CLK), .QN(n1096) );
  EDFFXL \targetY_reg[5][2]  ( .D(Y[2]), .E(n230), .CK(CLK), .QN(n1141) );
  EDFFXL \targetY_reg[5][0]  ( .D(Y[0]), .E(n230), .CK(CLK), .QN(n1084) );
  EDFFXL \targetY_reg[1][2]  ( .D(Y[2]), .E(n225), .CK(CLK), .QN(n1125) );
  EDFFXL \targetY_reg[1][0]  ( .D(Y[0]), .E(n225), .CK(CLK), .QN(n1088) );
  EDFFXL \targetX_reg[29][1]  ( .D(X[1]), .E(n233), .CK(CLK), .QN(n1101) );
  EDFFXL \targetX_reg[29][0]  ( .D(X[0]), .E(n233), .CK(CLK), .QN(n1076) );
  EDFFXL \targetX_reg[25][1]  ( .D(X[1]), .E(n228), .CK(CLK), .QN(n1161) );
  EDFFXL \targetX_reg[25][0]  ( .D(X[0]), .E(n228), .CK(CLK), .QN(n1080) );
  EDFFXL \targetX_reg[13][1]  ( .D(X[1]), .E(n231), .CK(CLK), .QN(n1185) );
  EDFFXL \targetX_reg[9][2]  ( .D(X[2]), .E(n226), .CK(CLK), .QN(n1205) );
  EDFFXL \targetX_reg[5][1]  ( .D(X[1]), .E(n230), .CK(CLK), .QN(n1189) );
  EDFFXL \targetX_reg[1][1]  ( .D(X[1]), .E(n225), .CK(CLK), .QN(n1117) );
  EDFFXL \targetX_reg[1][0]  ( .D(X[0]), .E(n225), .CK(CLK), .QN(n1113) );
  EDFFXL \targetY_reg[30][1]  ( .D(Y[1]), .E(n223), .CK(CLK), .QN(n1180) );
  EDFFXL \targetY_reg[22][2]  ( .D(Y[2]), .E(n222), .CK(CLK), .QN(n1144) );
  EDFFXL \targetY_reg[22][1]  ( .D(Y[1]), .E(n222), .CK(CLK), .QN(n1176) );
  EDFFXL \targetY_reg[20][2]  ( .D(Y[2]), .E(n217), .CK(CLK), .QN(n1143) );
  EDFFXL \targetY_reg[20][1]  ( .D(Y[1]), .E(n217), .CK(CLK), .QN(n1175) );
  EDFFXL \targetY_reg[14][2]  ( .D(Y[2]), .E(n221), .CK(CLK), .QN(n1104) );
  EDFFXL \targetY_reg[14][1]  ( .D(Y[1]), .E(n221), .CK(CLK), .QN(n1172) );
  EDFFXL \targetY_reg[14][0]  ( .D(Y[0]), .E(n221), .CK(CLK), .QN(n1091) );
  EDFFXL \targetY_reg[12][2]  ( .D(Y[2]), .E(n216), .CK(CLK), .QN(n1103) );
  EDFFXL \targetY_reg[12][1]  ( .D(Y[1]), .E(n216), .CK(CLK), .QN(n1171) );
  EDFFXL \targetY_reg[12][0]  ( .D(Y[0]), .E(n216), .CK(CLK), .QN(n1090) );
  EDFFXL \targetY_reg[4][2]  ( .D(Y[2]), .E(n215), .CK(CLK), .QN(n1139) );
  EDFFXL \targetY_reg[4][0]  ( .D(Y[0]), .E(n215), .CK(CLK), .QN(n1082) );
  EDFFXL \targetX_reg[30][1]  ( .D(X[1]), .E(n223), .CK(CLK), .QN(n1100) );
  EDFFXL \targetX_reg[30][0]  ( .D(X[0]), .E(n223), .CK(CLK), .QN(n1075) );
  EDFFXL \targetX_reg[22][1]  ( .D(X[1]), .E(n222), .CK(CLK), .QN(n1136) );
  EDFFXL \targetX_reg[22][0]  ( .D(X[0]), .E(n222), .CK(CLK), .QN(n1067) );
  EDFFXL \targetX_reg[20][1]  ( .D(X[1]), .E(n217), .CK(CLK), .QN(n1135) );
  EDFFXL \targetX_reg[20][0]  ( .D(X[0]), .E(n217), .CK(CLK), .QN(n1066) );
  EDFFXL \targetX_reg[14][1]  ( .D(X[1]), .E(n221), .CK(CLK), .QN(n1184) );
  EDFFXL \targetX_reg[12][1]  ( .D(X[1]), .E(n216), .CK(CLK), .QN(n1183) );
  EDFFXL \targetX_reg[4][1]  ( .D(X[1]), .E(n215), .CK(CLK), .QN(n1187) );
  EDFFXL \targetY_reg[3][2]  ( .D(Y[2]), .E(n235), .CK(CLK), .QN(n1126) );
  EDFFXL \targetY_reg[3][0]  ( .D(Y[0]), .E(n235), .CK(CLK), .QN(n1089) );
  EDFFXL \targetX_reg[27][1]  ( .D(X[1]), .E(n238), .CK(CLK), .QN(n1162) );
  EDFFXL \targetX_reg[27][0]  ( .D(X[0]), .E(n238), .CK(CLK), .QN(n1081) );
  EDFFXL \targetX_reg[19][1]  ( .D(X[1]), .E(n237), .CK(CLK), .QN(n1122) );
  EDFFXL \targetX_reg[19][0]  ( .D(X[0]), .E(n237), .CK(CLK), .QN(n1073) );
  EDFFXL \targetX_reg[3][1]  ( .D(X[1]), .E(n235), .CK(CLK), .QN(n1118) );
  EDFFXL \targetX_reg[3][0]  ( .D(X[0]), .E(n235), .CK(CLK), .QN(n1114) );
  EDFFXL \targetY_reg[10][2]  ( .D(Y[2]), .E(n211), .CK(CLK), .QN(n1164) );
  EDFFXL \targetY_reg[10][0]  ( .D(Y[0]), .E(n211), .CK(CLK), .QN(n1095) );
  EDFFXL \targetY_reg[8][2]  ( .D(Y[2]), .E(n206), .CK(CLK), .QN(n1163) );
  EDFFXL \targetY_reg[8][0]  ( .D(Y[0]), .E(n206), .CK(CLK), .QN(n1094) );
  EDFFXL \targetY_reg[0][2]  ( .D(Y[2]), .E(n205), .CK(CLK), .QN(n1123) );
  EDFFXL \targetY_reg[0][0]  ( .D(Y[0]), .E(n205), .CK(CLK), .QN(n1086) );
  EDFFXL \targetX_reg[26][1]  ( .D(X[1]), .E(n213), .CK(CLK), .QN(n1160) );
  EDFFXL \targetX_reg[26][0]  ( .D(X[0]), .E(n213), .CK(CLK), .QN(n1079) );
  EDFFXL \targetX_reg[18][1]  ( .D(X[1]), .E(n212), .CK(CLK), .QN(n1120) );
  EDFFXL \targetX_reg[18][0]  ( .D(X[0]), .E(n212), .CK(CLK), .QN(n1071) );
  EDFFXL \targetX_reg[16][1]  ( .D(X[1]), .E(n207), .CK(CLK), .QN(n1119) );
  EDFFXL \targetX_reg[16][0]  ( .D(X[0]), .E(n207), .CK(CLK), .QN(n1070) );
  EDFFXL \targetX_reg[10][1]  ( .D(X[1]), .E(n211), .CK(CLK), .QN(n1192) );
  EDFFXL \targetX_reg[8][1]  ( .D(X[1]), .E(n206), .CK(CLK), .QN(n1191) );
  EDFFXL \targetX_reg[0][1]  ( .D(X[1]), .E(n205), .CK(CLK), .QN(n1115) );
  EDFFXL \targetX_reg[0][0]  ( .D(X[0]), .E(n205), .CK(CLK), .QN(n1111) );
  EDFFXL \targetY_reg[15][1]  ( .D(Y[1]), .E(n241), .CK(CLK), .QN(n1174) );
  EDFFXL \targetX_reg[21][0]  ( .D(X[0]), .E(n232), .CK(CLK), .QN(n1068) );
  EDFFXL \targetX_reg[28][0]  ( .D(X[0]), .E(n218), .CK(CLK), .QN(n1074) );
  EDFFXL \targetY_reg[39][3]  ( .D(Y[3]), .E(n244), .CK(CLK), .Q(
        \targetY[39][3] ) );
  EDFFXL \targetY_reg[39][2]  ( .D(Y[2]), .E(n244), .CK(CLK), .Q(
        \targetY[39][2] ) );
  EDFFXL \targetY_reg[39][1]  ( .D(Y[1]), .E(n244), .CK(CLK), .Q(
        \targetY[39][1] ) );
  EDFFXL \targetY_reg[39][0]  ( .D(Y[0]), .E(n244), .CK(CLK), .Q(
        \targetY[39][0] ) );
  EDFFXL \targetX_reg[39][3]  ( .D(X[3]), .E(n244), .CK(CLK), .Q(
        \targetX[39][3] ) );
  EDFFXL \targetX_reg[39][2]  ( .D(X[2]), .E(n244), .CK(CLK), .Q(
        \targetX[39][2] ) );
  EDFFXL \targetX_reg[39][1]  ( .D(X[1]), .E(n244), .CK(CLK), .Q(
        \targetX[39][1] ) );
  EDFFXL \targetX_reg[39][0]  ( .D(X[0]), .E(n244), .CK(CLK), .Q(
        \targetX[39][0] ) );
  EDFFXL \targetY_reg[35][3]  ( .D(Y[3]), .E(n239), .CK(CLK), .Q(
        \targetY[35][3] ) );
  EDFFXL \targetY_reg[35][2]  ( .D(Y[2]), .E(n239), .CK(CLK), .Q(
        \targetY[35][2] ) );
  EDFFXL \targetY_reg[35][1]  ( .D(Y[1]), .E(n239), .CK(CLK), .Q(
        \targetY[35][1] ) );
  EDFFXL \targetY_reg[35][0]  ( .D(Y[0]), .E(n239), .CK(CLK), .Q(
        \targetY[35][0] ) );
  EDFFXL \targetX_reg[35][3]  ( .D(X[3]), .E(n239), .CK(CLK), .Q(
        \targetX[35][3] ) );
  EDFFXL \targetX_reg[35][2]  ( .D(X[2]), .E(n239), .CK(CLK), .Q(
        \targetX[35][2] ) );
  EDFFXL \targetX_reg[35][1]  ( .D(X[1]), .E(n239), .CK(CLK), .Q(
        \targetX[35][1] ) );
  EDFFXL \targetX_reg[35][0]  ( .D(X[0]), .E(n239), .CK(CLK), .Q(
        \targetX[35][0] ) );
  EDFFXL \targetY_reg[33][3]  ( .D(Y[3]), .E(n229), .CK(CLK), .Q(
        \targetY[33][3] ) );
  EDFFXL \targetX_reg[33][3]  ( .D(X[3]), .E(n229), .CK(CLK), .Q(
        \targetX[33][3] ) );
  EDFFXL \targetX_reg[33][2]  ( .D(X[2]), .E(n229), .CK(CLK), .Q(
        \targetX[33][2] ) );
  EDFFXL \targetY_reg[37][3]  ( .D(Y[3]), .E(n234), .CK(CLK), .Q(
        \targetY[37][3] ) );
  EDFFXL \targetX_reg[37][3]  ( .D(X[3]), .E(n234), .CK(CLK), .Q(
        \targetX[37][3] ) );
  EDFFXL \targetX_reg[37][2]  ( .D(X[2]), .E(n234), .CK(CLK), .Q(
        \targetX[37][2] ) );
  EDFFXL \targetY_reg[38][3]  ( .D(Y[3]), .E(n224), .CK(CLK), .Q(
        \targetY[38][3] ) );
  EDFFXL \targetX_reg[38][3]  ( .D(X[3]), .E(n224), .CK(CLK), .Q(
        \targetX[38][3] ) );
  EDFFXL \targetX_reg[38][2]  ( .D(X[2]), .E(n224), .CK(CLK), .Q(
        \targetX[38][2] ) );
  EDFFXL \targetY_reg[36][3]  ( .D(Y[3]), .E(n219), .CK(CLK), .Q(
        \targetY[36][3] ) );
  EDFFXL \targetX_reg[36][3]  ( .D(X[3]), .E(n219), .CK(CLK), .Q(
        \targetX[36][3] ) );
  EDFFXL \targetX_reg[36][2]  ( .D(X[2]), .E(n219), .CK(CLK), .Q(
        \targetX[36][2] ) );
  EDFFXL \targetY_reg[34][3]  ( .D(Y[3]), .E(n214), .CK(CLK), .Q(
        \targetY[34][3] ) );
  EDFFXL \targetY_reg[32][3]  ( .D(Y[3]), .E(n209), .CK(CLK), .Q(
        \targetY[32][3] ) );
  EDFFXL \targetX_reg[34][3]  ( .D(X[3]), .E(n214), .CK(CLK), .Q(
        \targetX[34][3] ) );
  EDFFXL \targetX_reg[34][0]  ( .D(X[0]), .E(n214), .CK(CLK), .Q(
        \targetX[34][0] ) );
  EDFFXL \targetX_reg[32][3]  ( .D(X[3]), .E(n209), .CK(CLK), .Q(
        \targetX[32][3] ) );
  EDFFXL \targetX_reg[32][2]  ( .D(X[2]), .E(n209), .CK(CLK), .Q(
        \targetX[32][2] ) );
  EDFFXL \targetX_reg[15][3]  ( .D(X[3]), .E(n241), .CK(CLK), .Q(
        \targetX[15][3] ) );
  EDFFXL \targetX_reg[7][3]  ( .D(X[3]), .E(n240), .CK(CLK), .Q(
        \targetX[7][3] ) );
  EDFFXL \targetY_reg[17][2]  ( .D(Y[2]), .E(n227), .CK(CLK), .Q(
        \targetY[17][2] ) );
  EDFFXL \targetY_reg[17][1]  ( .D(Y[1]), .E(n227), .CK(CLK), .Q(
        \targetY[17][1] ) );
  EDFFXL \targetY_reg[17][0]  ( .D(Y[0]), .E(n227), .CK(CLK), .Q(
        \targetY[17][0] ) );
  EDFFXL \targetY_reg[11][1]  ( .D(Y[1]), .E(n236), .CK(CLK), .Q(
        \targetY[11][1] ) );
  EDFFXL \targetX_reg[11][3]  ( .D(X[3]), .E(n236), .CK(CLK), .Q(
        \targetX[11][3] ) );
  EDFFXL \targetX_reg[11][0]  ( .D(X[0]), .E(n236), .CK(CLK), .Q(
        \targetX[11][0] ) );
  EDFFXL \targetY_reg[24][2]  ( .D(Y[2]), .E(n208), .CK(CLK), .Q(
        \targetY[24][2] ) );
  EDFFXL \targetY_reg[24][1]  ( .D(Y[1]), .E(n208), .CK(CLK), .Q(
        \targetY[24][1] ) );
  EDFFXL \targetY_reg[24][0]  ( .D(Y[0]), .E(n208), .CK(CLK), .Q(
        \targetY[24][0] ) );
  EDFFXL \targetY_reg[2][1]  ( .D(Y[1]), .E(n210), .CK(CLK), .Q(
        \targetY[2][1] ) );
  EDFFXL \targetY_reg[21][0]  ( .D(Y[0]), .E(n232), .CK(CLK), .Q(
        \targetY[21][0] ) );
  EDFFXL \targetY_reg[6][1]  ( .D(Y[1]), .E(n220), .CK(CLK), .Q(
        \targetY[6][1] ) );
  EDFFXL \targetX_reg[6][3]  ( .D(X[3]), .E(n220), .CK(CLK), .Q(
        \targetX[6][3] ) );
  EDFFXL \targetY_reg[28][2]  ( .D(Y[2]), .E(n218), .CK(CLK), .Q(
        \targetY[28][2] ) );
  EDFFXL \targetY_reg[28][0]  ( .D(Y[0]), .E(n218), .CK(CLK), .Q(
        \targetY[28][0] ) );
  EDFFXL \targetX_reg[13][3]  ( .D(X[3]), .E(n231), .CK(CLK), .Q(
        \targetX[13][3] ) );
  EDFFXL \targetX_reg[9][3]  ( .D(X[3]), .E(n226), .CK(CLK), .Q(
        \targetX[9][3] ) );
  EDFFXL \targetX_reg[5][3]  ( .D(X[3]), .E(n230), .CK(CLK), .Q(
        \targetX[5][3] ) );
  EDFFXL \targetX_reg[14][3]  ( .D(X[3]), .E(n221), .CK(CLK), .Q(
        \targetX[14][3] ) );
  EDFFXL \targetX_reg[12][3]  ( .D(X[3]), .E(n216), .CK(CLK), .Q(
        \targetX[12][3] ) );
  EDFFXL \targetX_reg[4][3]  ( .D(X[3]), .E(n215), .CK(CLK), .Q(
        \targetX[4][3] ) );
  EDFFXL \targetX_reg[10][3]  ( .D(X[3]), .E(n211), .CK(CLK), .Q(
        \targetX[10][3] ) );
  EDFFXL \targetX_reg[8][3]  ( .D(X[3]), .E(n206), .CK(CLK), .Q(
        \targetX[8][3] ) );
  DFFRX1 optimise_reg ( .D(n245), .CK(CLK), .RN(n1568), .Q(optimise), .QN(
        n1509) );
  DFFRX1 \max_covered_1_reg[5]  ( .D(n302), .CK(CLK), .RN(n1568), .Q(n1512), 
        .QN(n187) );
  DFFRX1 \max_covered_1_reg[4]  ( .D(n303), .CK(CLK), .RN(n1568), .QN(n186) );
  DFFRX1 \max_covered_1_reg[3]  ( .D(n304), .CK(CLK), .RN(n1568), .Q(n1516), 
        .QN(n185) );
  DFFRX1 \max_covered_1_reg[2]  ( .D(n305), .CK(CLK), .RN(n1568), .QN(n263) );
  DFFRX1 \max_covered_1_reg[1]  ( .D(n306), .CK(CLK), .RN(n1568), .QN(n264) );
  DFFRX1 \max_covered_1_reg[0]  ( .D(n307), .CK(CLK), .RN(n1568), .QN(n265) );
  DFFRX1 \max_covered_2_reg[5]  ( .D(n278), .CK(CLK), .RN(n1568), .Q(n1500), 
        .QN(n202) );
  DFFRX1 \max_covered_2_reg[4]  ( .D(n279), .CK(CLK), .RN(n1568), .QN(n201) );
  DFFRX1 \max_covered_2_reg[3]  ( .D(n280), .CK(CLK), .RN(n1568), .QN(n200) );
  DFFRX1 \max_covered_2_reg[2]  ( .D(n281), .CK(CLK), .RN(n1568), .QN(n199) );
  DFFRX1 \max_covered_2_reg[1]  ( .D(n282), .CK(CLK), .RN(n1568), .QN(n198) );
  DFFRX1 \max_covered_2_reg[0]  ( .D(n283), .CK(CLK), .RN(n1568), .QN(n197) );
  DFFRX1 \yMax2_reg[3]  ( .D(n318), .CK(CLK), .RN(n1568), .QN(n1555) );
  DFFRX1 \yMax2_reg[2]  ( .D(n308), .CK(CLK), .RN(n1568), .QN(n1553) );
  DFFRX1 \yMax2_reg[0]  ( .D(n312), .CK(CLK), .RN(n1568), .QN(n1554) );
  DFFRX1 \yMax1_reg[3]  ( .D(n300), .CK(CLK), .RN(n1568), .QN(n1560) );
  DFFRX1 \yMax1_reg[2]  ( .D(n286), .CK(CLK), .RN(n1568), .QN(n1565) );
  DFFRX1 \yMax1_reg[0]  ( .D(n290), .CK(CLK), .RN(n1568), .QN(n1566) );
  DFFRX1 \xMax2_reg[3]  ( .D(n277), .CK(CLK), .RN(n1568), .QN(n1556) );
  DFFRX1 \xMax2_reg[2]  ( .D(n284), .CK(CLK), .RN(n1568), .QN(n1557) );
  DFFRX1 \xMax2_reg[1]  ( .D(n315), .CK(CLK), .RN(n1568), .QN(n1558) );
  DFFRX1 \xMax2_reg[0]  ( .D(n319), .CK(CLK), .RN(n1568), .QN(n1559) );
  DFFRX1 \xMax1_reg[3]  ( .D(n297), .CK(CLK), .RN(n1568), .QN(n1564) );
  DFFRX1 \xMax1_reg[2]  ( .D(n285), .CK(CLK), .RN(n1568), .QN(n1561) );
  DFFRX1 \xMax1_reg[1]  ( .D(n293), .CK(CLK), .RN(n1568), .QN(n1562) );
  DFFRX1 \xMax1_reg[0]  ( .D(n295), .CK(CLK), .RN(n1568), .QN(n1563) );
  DFFRX1 \count_reg[3]  ( .D(n328), .CK(CLK), .RN(n1379), .Q(count[3]), .QN(
        n259) );
  DFFRX1 \state_reg[2]  ( .D(nextState[2]), .CK(CLK), .RN(n1378), .Q(state[2]), 
        .QN(n1045) );
  DFFRX2 \count_reg[4]  ( .D(n327), .CK(CLK), .RN(n1379), .Q(count[4]), .QN(
        n258) );
  DFFRX2 \count_reg[2]  ( .D(n329), .CK(CLK), .RN(n1379), .Q(count[2]), .QN(
        n260) );
  DFFRX2 \count_reg[5]  ( .D(n326), .CK(CLK), .RN(n1379), .Q(count[5]), .QN(
        n257) );
  ADDFHX2 \r399/U2_3  ( .A(n1571), .B(n1385), .CI(\r399/carry[3] ), .CO(
        \r399/carry[4] ), .S(N829) );
  ADDFHX4 \r401/U2_3  ( .A(n1575), .B(n1040), .CI(\r401/carry[3] ), .CO(
        \r401/carry[4] ), .S(N846) );
  ADDFHX4 \r404/U2_2  ( .A(C2X[2]), .B(n1041), .CI(\r404/carry[2] ), .CO(
        \r404/carry[3] ), .S(N950) );
  ADDFHX4 \r399/U2_2  ( .A(C1X[2]), .B(n1041), .CI(\r399/carry[2] ), .CO(
        \r399/carry[3] ), .S(N828) );
  ADDFX2 \r401/U2_0  ( .A(n1578), .B(n1360), .CI(1'b1), .CO(\r401/carry[1] ), 
        .S(N843) );
  MXI2X1 U970 ( .A(n1276), .B(n1281), .S0(n258), .Y(n1063) );
  MX4X1 U971 ( .A(n1275), .B(n1273), .C(n1274), .D(n1272), .S0(n1377), .S1(
        n1362), .Y(n1276) );
  MXI3X2 U972 ( .A(n1341), .B(n1346), .C(n1334), .S0(n258), .S1(count[5]), .Y(
        n1041) );
  MXI3X2 U973 ( .A(n1302), .B(n1307), .C(n1295), .S0(n258), .S1(count[5]), .Y(
        n1040) );
  BUFX20 U974 ( .A(n1364), .Y(n1039) );
  CLKBUFX2 U975 ( .A(n1061), .Y(n1364) );
  MXI4X1 U976 ( .A(n1111), .B(n1112), .C(n1113), .D(n1114), .S0(n1367), .S1(
        n1372), .Y(n1319) );
  NAND2X1 U977 ( .A(n1252), .B(n1253), .Y(\r406/carry[1] ) );
  INVX1 U978 ( .A(n1360), .Y(n1252) );
  MX4XL U979 ( .A(\targetY[24][0] ), .B(\targetY[26][0] ), .C(\targetY[25][0] ), .D(\targetY[27][0] ), .S0(n1368), .S1(n1251), .Y(n1261) );
  MX4XL U980 ( .A(\targetY[16][0] ), .B(\targetY[18][0] ), .C(\targetY[17][0] ), .D(\targetY[19][0] ), .S0(n1368), .S1(n1375), .Y(n1263) );
  MX4X1 U981 ( .A(\targetY[8][1] ), .B(\targetY[10][1] ), .C(\targetY[9][1] ), 
        .D(\targetY[11][1] ), .S0(n1366), .S1(n1374), .Y(n1278) );
  MX3X2 U982 ( .A(n1328), .B(n1333), .C(n1321), .S0(n258), .S1(count[5]), .Y(
        n1098) );
  MX4X2 U983 ( .A(n1319), .B(n1317), .C(n1318), .D(n1316), .S0(n1377), .S1(
        n1363), .Y(n1320) );
  MX4X1 U984 ( .A(n1263), .B(n1261), .C(n1262), .D(n1260), .S0(n1377), .S1(
        n1362), .Y(n1264) );
  MX4X1 U985 ( .A(n1268), .B(n1266), .C(n1267), .D(n1265), .S0(n1377), .S1(
        n1362), .Y(n1269) );
  BUFX2 U986 ( .A(count[0]), .Y(n1376) );
  XNOR2X2 U987 ( .A(n1387), .B(n1582), .Y(N948) );
  XNOR2X2 U988 ( .A(n1383), .B(n1574), .Y(N826) );
  CLKINVX1 U989 ( .A(n1586), .Y(n1253) );
  OAI31X1 U990 ( .A0(n1448), .A1(n1433), .A2(n1405), .B0(n1439), .Y(n1418) );
  BUFX4 U991 ( .A(n1061), .Y(n1365) );
  CLKBUFX8 U992 ( .A(n1365), .Y(n1368) );
  BUFX4 U993 ( .A(n1376), .Y(n1375) );
  BUFX12 U994 ( .A(n1365), .Y(n1367) );
  BUFX4 U995 ( .A(n1365), .Y(n1366) );
  MXI3X2 U996 ( .A(n1289), .B(n1294), .C(n1282), .S0(n258), .S1(count[5]), .Y(
        n1042) );
  BUFX4 U997 ( .A(n1376), .Y(n1374) );
  MX3X1 U998 ( .A(n1354), .B(n1359), .C(n1347), .S0(n258), .S1(count[5]), .Y(
        n1065) );
  CLKMX2X2 U999 ( .A(n1270), .B(n1271), .S0(n1363), .Y(n1043) );
  MXI2X2 U1000 ( .A(n1063), .B(n1043), .S0(count[5]), .Y(n1064) );
  CLKINVX1 U1001 ( .A(count[0]), .Y(n1382) );
  CLKINVX1 U1002 ( .A(n262), .Y(n1251) );
  CLKBUFX6 U1003 ( .A(count[3]), .Y(n1377) );
  BUFX16 U1004 ( .A(n1580), .Y(C2X[2]) );
  BUFX16 U1005 ( .A(n1584), .Y(C2Y[2]) );
  BUFX16 U1006 ( .A(n1585), .Y(C2Y[1]) );
  BUFX16 U1007 ( .A(n1573), .Y(C1X[1]) );
  BUFX16 U1008 ( .A(n1572), .Y(C1X[2]) );
  AND2X2 U1009 ( .A(n1520), .B(n1521), .Y(n244) );
  INVX6 U1010 ( .A(RST), .Y(n1568) );
  CLKBUFX3 U1011 ( .A(n1062), .Y(n1047) );
  INVXL U1012 ( .A(n1061), .Y(n1062) );
  INVX2 U1013 ( .A(n1064), .Y(n1389) );
  NOR2X2 U1014 ( .A(n1528), .B(n1532), .Y(n219) );
  NOR2X2 U1015 ( .A(n1523), .B(n1527), .Y(n238) );
  NOR2X2 U1016 ( .A(n1524), .B(n1531), .Y(n222) );
  NOR2X2 U1017 ( .A(n1525), .B(n1529), .Y(n231) );
  NOR2X2 U1018 ( .A(n1522), .B(n1526), .Y(n240) );
  NOR2X2 U1019 ( .A(n1528), .B(n1533), .Y(n214) );
  NOR2X2 U1020 ( .A(n1523), .B(n1529), .Y(n233) );
  NOR2X2 U1021 ( .A(n1522), .B(n1524), .Y(n242) );
  NOR2X2 U1022 ( .A(n1525), .B(n1530), .Y(n226) );
  NOR2X2 U1023 ( .A(n1526), .B(n1527), .Y(n235) );
  NOR2X2 U1024 ( .A(n1528), .B(n1534), .Y(n209) );
  NOR2X2 U1025 ( .A(n1523), .B(n1533), .Y(n213) );
  NOR2X2 U1026 ( .A(n1524), .B(n1527), .Y(n237) );
  NOR2X2 U1027 ( .A(n1526), .B(n1529), .Y(n230) );
  NOR2X2 U1028 ( .A(n1525), .B(n1531), .Y(n221) );
  NOR2X2 U1029 ( .A(n1528), .B(n1529), .Y(n234) );
  NOR2X2 U1030 ( .A(n1522), .B(n1523), .Y(n243) );
  NOR2X2 U1031 ( .A(n1524), .B(n1534), .Y(n207) );
  NOR2X2 U1032 ( .A(n1526), .B(n1530), .Y(n225) );
  NOR2X2 U1033 ( .A(n1525), .B(n1532), .Y(n216) );
  NOR4X2 U1034 ( .A(n1377), .B(count[4]), .C(n1522), .D(n257), .Y(n1521) );
  OAI21X1 U1035 ( .A0(n1481), .A1(n1437), .B0(n1480), .Y(n1464) );
  NOR2X2 U1036 ( .A(n1528), .B(n1531), .Y(n224) );
  NOR2X2 U1037 ( .A(n1523), .B(n1530), .Y(n228) );
  NOR2X2 U1038 ( .A(n1524), .B(n1533), .Y(n212) );
  NOR2X2 U1039 ( .A(n1526), .B(n1532), .Y(n215) );
  NOR2X2 U1040 ( .A(n1525), .B(n1534), .Y(n206) );
  NOR3X2 U1041 ( .A(n1396), .B(n1430), .C(n1431), .Y(n1397) );
  NAND3X2 U1042 ( .A(n1415), .B(n1497), .C(optimise), .Y(n1496) );
  NAND3X2 U1043 ( .A(n1508), .B(n1509), .C(n1415), .Y(n1450) );
  NOR3X2 U1044 ( .A(state[0]), .B(state[1]), .C(n1045), .Y(n1415) );
  BUFX12 U1045 ( .A(n1587), .Y(DONE) );
  OAI21X1 U1046 ( .A0(n1492), .A1(n1437), .B0(n1485), .Y(n1458) );
  NOR2X2 U1047 ( .A(n1528), .B(n1530), .Y(n229) );
  NOR2X2 U1048 ( .A(n1527), .B(n1528), .Y(n239) );
  NAND4BX2 U1049 ( .AN(n257), .B(n1520), .C(n259), .D(n258), .Y(n1528) );
  NOR2X2 U1050 ( .A(n1523), .B(n1531), .Y(n223) );
  NOR2X2 U1051 ( .A(n1524), .B(n1532), .Y(n217) );
  NOR2X2 U1052 ( .A(n1525), .B(n1533), .Y(n211) );
  NOR2X2 U1053 ( .A(n1526), .B(n1534), .Y(n205) );
  OA21X2 U1054 ( .A0(n1494), .A1(n1495), .B0(n1567), .Y(n1456) );
  OAI21X1 U1055 ( .A0(n1434), .A1(n1410), .B0(n1411), .Y(n1439) );
  NOR3X2 U1056 ( .A(n1472), .B(n1481), .C(n1410), .Y(n1468) );
  INVX3 U1057 ( .A(n1433), .Y(n1410) );
  BUFX12 U1058 ( .A(n1578), .Y(C1Y[0]) );
  BUFX12 U1059 ( .A(n1577), .Y(C1Y[1]) );
  INVX16 U1060 ( .A(n204), .Y(C2X[3]) );
  INVX12 U1061 ( .A(n247), .Y(C2Y[3]) );
  INVX12 U1062 ( .A(n270), .Y(C1Y[3]) );
  INVX12 U1063 ( .A(n266), .Y(C1X[3]) );
  BUFX12 U1064 ( .A(n1576), .Y(C1Y[2]) );
  BUFX12 U1065 ( .A(n1581), .Y(C2X[1]) );
  NOR2X2 U1066 ( .A(n1523), .B(n1532), .Y(n218) );
  NOR2X2 U1067 ( .A(n1523), .B(n1534), .Y(n208) );
  NAND3X2 U1068 ( .A(count[4]), .B(n1377), .C(n1535), .Y(n1523) );
  NOR2X2 U1069 ( .A(n1524), .B(n1529), .Y(n232) );
  NOR2X2 U1070 ( .A(n1524), .B(n1530), .Y(n227) );
  NAND3X2 U1071 ( .A(n259), .B(count[4]), .C(n1535), .Y(n1524) );
  NOR2X2 U1072 ( .A(n1522), .B(n1525), .Y(n241) );
  NOR2X2 U1073 ( .A(n1525), .B(n1527), .Y(n236) );
  NAND3X2 U1074 ( .A(n258), .B(n1377), .C(n1535), .Y(n1525) );
  NOR2X2 U1075 ( .A(n1526), .B(n1531), .Y(n220) );
  NOR2X2 U1076 ( .A(n1526), .B(n1533), .Y(n210) );
  NAND3X2 U1077 ( .A(n259), .B(n258), .C(n1535), .Y(n1526) );
  INVX12 U1078 ( .A(n1253), .Y(C2Y[0]) );
  OAI31X1 U1079 ( .A0(n1405), .A1(n1430), .A2(n1433), .B0(n1432), .Y(n1394) );
  NOR3X2 U1080 ( .A(state[1]), .B(state[2]), .C(state[0]), .Y(n1405) );
  OA21X2 U1081 ( .A0(n1494), .A1(n1495), .B0(n1455), .Y(n1417) );
  INVX12 U1082 ( .A(n1255), .Y(C2X[0]) );
  CLKINVX1 U1083 ( .A(n1582), .Y(n1255) );
  INVX12 U1084 ( .A(n1256), .Y(C1X[0]) );
  CLKINVX1 U1085 ( .A(n1574), .Y(n1256) );
  BUFX12 U1086 ( .A(n1376), .Y(n1369) );
  MXI4X2 U1087 ( .A(n1066), .B(n1067), .C(n1068), .D(n1069), .S0(n1367), .S1(
        n1373), .Y(n1313) );
  MXI4X2 U1088 ( .A(n1074), .B(n1075), .C(n1076), .D(n1077), .S0(n1367), .S1(
        n1373), .Y(n1311) );
  MXI4X2 U1089 ( .A(n1078), .B(n1079), .C(n1080), .D(n1081), .S0(n1367), .S1(
        n1373), .Y(n1312) );
  BUFX20 U1090 ( .A(n1369), .Y(n1373) );
  NOR2X2 U1091 ( .A(N982), .B(N983), .Y(n1416) );
  OAI32X2 U1092 ( .A0(n1391), .A1(len1[0]), .A2(n1390), .B0(len1[4]), .B1(
        n1390), .Y(N982) );
  BUFX12 U1093 ( .A(n1370), .Y(n1371) );
  AOI31XL U1094 ( .A0(state[0]), .A1(n1046), .A2(state[2]), .B0(n1405), .Y(
        n1404) );
  BUFX12 U1095 ( .A(n1369), .Y(n1372) );
  MX4X1 U1096 ( .A(n1280), .B(n1278), .C(n1279), .D(n1277), .S0(n1377), .S1(
        n1362), .Y(n1281) );
  INVXL U1097 ( .A(n1397), .Y(n1401) );
  INVXL U1098 ( .A(n1468), .Y(n1475) );
  NAND2XL U1099 ( .A(n1483), .B(n1410), .Y(n1485) );
  INVXL U1100 ( .A(n1450), .Y(n1494) );
  INVXL U1101 ( .A(n1496), .Y(n1495) );
  AOI2BB1XL U1102 ( .A0N(n1431), .A1N(n1452), .B0(n1405), .Y(n1483) );
  INVX1 U1103 ( .A(n1415), .Y(n1412) );
  INVXL U1104 ( .A(n1521), .Y(n1409) );
  MXI2XL U1105 ( .A(n1452), .B(n1453), .S0(n1410), .Y(n1451) );
  NAND3XL U1106 ( .A(n1539), .B(n1540), .C(n1521), .Y(n1538) );
  MXI2X2 U1107 ( .A(n1309), .B(n1310), .S0(n1363), .Y(n1308) );
  MXI2X1 U1108 ( .A(n1258), .B(n1259), .S0(n1363), .Y(n1257) );
  MXI4XL U1109 ( .A(n1099), .B(n1100), .C(n1101), .D(n1102), .S0(n1367), .S1(
        n1372), .Y(n1324) );
  INVX1 U1110 ( .A(n1098), .Y(n1384) );
  MXI4XL U1111 ( .A(n1107), .B(n1108), .C(n1109), .D(n1110), .S0(n1039), .S1(
        n1372), .Y(n1337) );
  MXI4XL U1112 ( .A(n1131), .B(n1132), .C(n1133), .D(n1134), .S0(n1039), .S1(
        n1369), .Y(n1350) );
  MXI4XL U1113 ( .A(n1151), .B(n1152), .C(n1153), .D(n1154), .S0(n1039), .S1(
        n1369), .Y(n1345) );
  MXI2XL U1114 ( .A(n1553), .B(n248), .S0(n1417), .Y(n308) );
  MXI2XL U1115 ( .A(n1441), .B(n249), .S0(n1417), .Y(n310) );
  MXI2XL U1116 ( .A(n1554), .B(n250), .S0(n1417), .Y(n312) );
  MXI2XL U1117 ( .A(n1555), .B(n247), .S0(n1417), .Y(n318) );
  MXI2XL U1118 ( .A(n1556), .B(n204), .S0(n1417), .Y(n277) );
  MXI2XL U1119 ( .A(n1557), .B(n274), .S0(n1417), .Y(n284) );
  MXI2XL U1120 ( .A(n1558), .B(n275), .S0(n1417), .Y(n315) );
  MXI2XL U1121 ( .A(n1559), .B(n276), .S0(n1417), .Y(n319) );
  MXI2XL U1122 ( .A(n1560), .B(n270), .S0(n1456), .Y(n300) );
  MXI2XL U1123 ( .A(n1561), .B(n267), .S0(n1456), .Y(n285) );
  MXI2XL U1124 ( .A(n1562), .B(n268), .S0(n1456), .Y(n293) );
  MXI2XL U1125 ( .A(n1563), .B(n269), .S0(n1456), .Y(n295) );
  MXI2XL U1126 ( .A(n1564), .B(n266), .S0(n1456), .Y(n297) );
  MXI2XL U1127 ( .A(n1565), .B(n271), .S0(n1456), .Y(n286) );
  MXI2XL U1128 ( .A(n1487), .B(n272), .S0(n1456), .Y(n288) );
  MXI2XL U1129 ( .A(n1566), .B(n273), .S0(n1456), .Y(n290) );
  AO21XL U1130 ( .A0(n275), .A1(n1397), .B0(n1402), .Y(n1428) );
  AO21XL U1131 ( .A0(n276), .A1(n1397), .B0(n1396), .Y(n1402) );
  OAI211XL U1132 ( .A0(n1556), .A1(n1394), .B0(n1398), .C0(n1399), .Y(n333) );
  MXI2XL U1133 ( .A(n1396), .B(n1397), .S0(n276), .Y(n1395) );
  OAI211XL U1134 ( .A0(n1564), .A1(n1464), .B0(n1465), .C0(n1466), .Y(n298) );
  NAND3BXL U1135 ( .AN(n267), .B(n1467), .C(n1468), .Y(n1466) );
  OAI2BB1XL U1136 ( .A0N(n1468), .A1N(n269), .B0(n1480), .Y(n1469) );
  MXI2XL U1137 ( .A(n1472), .B(n1468), .S0(n269), .Y(n1471) );
  AO21XL U1138 ( .A0(n1468), .A1(n268), .B0(n1469), .Y(n1477) );
  MX2XL U1139 ( .A(n1439), .B(n1440), .S0(n250), .Y(n1438) );
  MXI2XL U1140 ( .A(n255), .B(n198), .S0(n1496), .Y(n282) );
  MXI2XL U1141 ( .A(n254), .B(n199), .S0(n1496), .Y(n281) );
  MXI2XL U1142 ( .A(n253), .B(n200), .S0(n1496), .Y(n280) );
  MXI2XL U1143 ( .A(n252), .B(n201), .S0(n1496), .Y(n279) );
  MXI2XL U1144 ( .A(n256), .B(n197), .S0(n1496), .Y(n283) );
  OAI211XL U1145 ( .A0(n1555), .A1(n1418), .B0(n1419), .C0(n1420), .Y(n317) );
  OAI2BB1XL U1146 ( .A0N(n1422), .A1N(n250), .B0(n1439), .Y(n1443) );
  MXI2XL U1147 ( .A(n252), .B(n186), .S0(n1450), .Y(n303) );
  MXI2XL U1148 ( .A(n253), .B(n185), .S0(n1450), .Y(n304) );
  MXI2XL U1149 ( .A(n254), .B(n263), .S0(n1450), .Y(n305) );
  MXI2XL U1150 ( .A(n255), .B(n264), .S0(n1450), .Y(n306) );
  MXI2XL U1151 ( .A(n256), .B(n265), .S0(n1450), .Y(n307) );
  AOI31XL U1152 ( .A0(n1542), .A1(n1539), .A2(n1415), .B0(n1405), .Y(n1541) );
  NAND3XL U1153 ( .A(state[0]), .B(n1045), .C(n1521), .Y(n1537) );
  NAND2BX4 U1154 ( .AN(n1383), .B(n1256), .Y(\r399/carry[1] ) );
  MXI4X1 U1155 ( .A(n1070), .B(n1071), .C(n1072), .D(n1073), .S0(n1367), .S1(
        n1251), .Y(n1314) );
  MXI4XL U1156 ( .A(n1082), .B(n1083), .C(n1084), .D(n1085), .S0(n1368), .S1(
        n1375), .Y(n1267) );
  MXI4XL U1157 ( .A(n1086), .B(n1087), .C(n1088), .D(n1089), .S0(n1368), .S1(
        n1375), .Y(n1268) );
  MXI4XL U1158 ( .A(n1090), .B(n1091), .C(n1092), .D(n1093), .S0(n1368), .S1(
        n1375), .Y(n1265) );
  MXI4XL U1159 ( .A(n1094), .B(n1095), .C(n1096), .D(n1097), .S0(n1368), .S1(
        n1375), .Y(n1266) );
  MXI4XL U1160 ( .A(n1103), .B(n1104), .C(n1105), .D(n1106), .S0(n1367), .S1(
        n1374), .Y(n1290) );
  MXI4XL U1161 ( .A(n1115), .B(n1116), .C(n1117), .D(n1118), .S0(n1367), .S1(
        n1372), .Y(n1332) );
  MXI4XL U1162 ( .A(n1119), .B(n1120), .C(n1121), .D(n1122), .S0(n1367), .S1(
        n1372), .Y(n1327) );
  MXI4XL U1163 ( .A(n1123), .B(n1124), .C(n1125), .D(n1126), .S0(n1367), .S1(
        n1374), .Y(n1293) );
  MXI4XL U1164 ( .A(n1127), .B(n1128), .C(n1129), .D(n1130), .S0(n1039), .S1(
        n1372), .Y(n1340) );
  MXI4XL U1165 ( .A(n1135), .B(n1136), .C(n1137), .D(n1138), .S0(n1367), .S1(
        n1372), .Y(n1326) );
  MXI4XL U1166 ( .A(n1139), .B(n1140), .C(n1141), .D(n1142), .S0(n1367), .S1(
        n1374), .Y(n1292) );
  MXI4XL U1167 ( .A(n1143), .B(n1144), .C(n1145), .D(n1146), .S0(n1366), .S1(
        n1374), .Y(n1287) );
  MXI4XL U1168 ( .A(n1147), .B(n1148), .C(n1149), .D(n1150), .S0(n1039), .S1(
        n1372), .Y(n1339) );
  MXI4XL U1169 ( .A(n1155), .B(n1156), .C(n1157), .D(n1158), .S0(n1039), .S1(
        n1369), .Y(n1352) );
  MXI4XL U1170 ( .A(n1159), .B(n1160), .C(n1161), .D(n1162), .S0(n1367), .S1(
        n1372), .Y(n1325) );
  MXI4XL U1171 ( .A(n1163), .B(n1164), .C(n1165), .D(n1166), .S0(n1367), .S1(
        n1374), .Y(n1291) );
  MXI4XL U1172 ( .A(n1167), .B(n1168), .C(n1169), .D(n1170), .S0(n1039), .S1(
        n1372), .Y(n1338) );
  MX4X1 U1173 ( .A(\targetY[28][0] ), .B(\targetY[30][0] ), .C(
        \targetY[29][0] ), .D(\targetY[31][0] ), .S0(n1368), .S1(n1251), .Y(
        n1260) );
  MXI4XL U1174 ( .A(n1171), .B(n1172), .C(n1173), .D(n1174), .S0(n1368), .S1(
        n1375), .Y(n1277) );
  MXI4XL U1175 ( .A(n1175), .B(n1176), .C(n1177), .D(n1178), .S0(n1368), .S1(
        n1375), .Y(n1274) );
  MXI4XL U1176 ( .A(\targetX[36][0] ), .B(\targetX[38][0] ), .C(
        \targetX[37][0] ), .D(\targetX[39][0] ), .S0(n1367), .S1(n1371), .Y(
        n1310) );
  MXI4XL U1177 ( .A(\targetX[36][1] ), .B(\targetX[38][1] ), .C(
        \targetX[37][1] ), .D(\targetX[39][1] ), .S0(n1367), .S1(n1371), .Y(
        n1323) );
  MXI4XL U1178 ( .A(\targetY[36][2] ), .B(\targetY[38][2] ), .C(
        \targetY[37][2] ), .D(\targetY[39][2] ), .S0(n1366), .S1(n1371), .Y(
        n1284) );
  MXI4XL U1179 ( .A(\targetX[36][2] ), .B(\targetX[38][2] ), .C(
        \targetX[37][2] ), .D(\targetX[39][2] ), .S0(n1039), .S1(n1371), .Y(
        n1336) );
  MXI4XL U1180 ( .A(\targetY[32][0] ), .B(\targetY[34][0] ), .C(
        \targetY[33][0] ), .D(\targetY[35][0] ), .S0(n1039), .S1(n1371), .Y(
        n1258) );
  MXI4XL U1181 ( .A(\targetX[32][0] ), .B(\targetX[34][0] ), .C(
        \targetX[33][0] ), .D(\targetX[35][0] ), .S0(n1367), .S1(n1371), .Y(
        n1309) );
  MXI4XL U1182 ( .A(\targetX[32][1] ), .B(\targetX[34][1] ), .C(
        \targetX[33][1] ), .D(\targetX[35][1] ), .S0(n1039), .S1(n1371), .Y(
        n1322) );
  MXI4XL U1183 ( .A(\targetY[32][2] ), .B(\targetY[34][2] ), .C(
        \targetY[33][2] ), .D(\targetY[35][2] ), .S0(n1366), .S1(n1371), .Y(
        n1283) );
  MXI4XL U1184 ( .A(\targetX[32][2] ), .B(\targetX[34][2] ), .C(
        \targetX[33][2] ), .D(\targetX[35][2] ), .S0(n1039), .S1(n1371), .Y(
        n1335) );
  MXI4XL U1185 ( .A(\targetY[36][0] ), .B(\targetY[38][0] ), .C(
        \targetY[37][0] ), .D(\targetY[39][0] ), .S0(n1039), .S1(n1369), .Y(
        n1259) );
  MXI4XL U1186 ( .A(n1179), .B(n1180), .C(n1181), .D(n1182), .S0(n1039), .S1(
        n1375), .Y(n1272) );
  MX4XL U1187 ( .A(\targetY[16][2] ), .B(\targetY[18][2] ), .C(
        \targetY[17][2] ), .D(\targetY[19][2] ), .S0(n1366), .S1(n1374), .Y(
        n1288) );
  MX4XL U1188 ( .A(\targetY[24][2] ), .B(\targetY[26][2] ), .C(
        \targetY[25][2] ), .D(\targetY[27][2] ), .S0(n1366), .S1(n1374), .Y(
        n1286) );
  MX4XL U1189 ( .A(\targetY[28][2] ), .B(\targetY[30][2] ), .C(
        \targetY[29][2] ), .D(\targetY[31][2] ), .S0(n1367), .S1(n1374), .Y(
        n1285) );
  MXI4XL U1190 ( .A(n1183), .B(n1184), .C(n1185), .D(n1186), .S0(n1367), .S1(
        n1372), .Y(n1329) );
  MXI4XL U1191 ( .A(n1187), .B(n1188), .C(n1189), .D(n1190), .S0(n1367), .S1(
        n1372), .Y(n1331) );
  MXI4XL U1192 ( .A(n1191), .B(n1192), .C(n1193), .D(n1194), .S0(n1367), .S1(
        n1372), .Y(n1330) );
  MXI4XL U1193 ( .A(n1195), .B(n1196), .C(n1197), .D(n1198), .S0(n1039), .S1(
        n1369), .Y(n1342) );
  MXI4XL U1194 ( .A(n1199), .B(n1200), .C(n1201), .D(n1202), .S0(n1039), .S1(
        n1369), .Y(n1344) );
  MXI4XL U1195 ( .A(n1203), .B(n1204), .C(n1205), .D(n1206), .S0(n1039), .S1(
        n1369), .Y(n1343) );
  MX4XL U1196 ( .A(\targetX[12][3] ), .B(\targetX[14][3] ), .C(
        \targetX[13][3] ), .D(\targetX[15][3] ), .S0(n1039), .S1(n1369), .Y(
        n1355) );
  MX4XL U1197 ( .A(\targetX[4][3] ), .B(\targetX[6][3] ), .C(\targetX[5][3] ), 
        .D(\targetX[7][3] ), .S0(n1039), .S1(n1369), .Y(n1357) );
  MX4XL U1198 ( .A(\targetX[8][3] ), .B(\targetX[10][3] ), .C(\targetX[9][3] ), 
        .D(\targetX[11][3] ), .S0(n1039), .S1(n1369), .Y(n1356) );
  CLKINVX4 U1199 ( .A(n1361), .Y(N903) );
  MXI4XL U1200 ( .A(n1207), .B(n1208), .C(n1209), .D(n1210), .S0(n1039), .S1(
        n1373), .Y(n1303) );
  MXI4XL U1201 ( .A(n1211), .B(n1212), .C(n1213), .D(n1214), .S0(n1367), .S1(
        n1373), .Y(n1301) );
  MXI4XL U1202 ( .A(n1215), .B(n1216), .C(n1217), .D(n1218), .S0(n1368), .S1(
        n1374), .Y(n1299) );
  MXI4XL U1203 ( .A(n1219), .B(n1220), .C(n1221), .D(n1222), .S0(n1367), .S1(
        n1374), .Y(n1298) );
  MXI4XL U1204 ( .A(n1223), .B(n1224), .C(n1225), .D(n1226), .S0(n1367), .S1(
        n1373), .Y(n1306) );
  MXI4XL U1205 ( .A(n1227), .B(n1228), .C(n1229), .D(n1230), .S0(n1039), .S1(
        n1373), .Y(n1305) );
  MXI4XL U1206 ( .A(n1231), .B(n1232), .C(n1233), .D(n1234), .S0(n1039), .S1(
        n1373), .Y(n1300) );
  MXI4XL U1207 ( .A(n1235), .B(n1236), .C(n1237), .D(n1238), .S0(n1039), .S1(
        n1375), .Y(n1358) );
  MXI4XL U1208 ( .A(n1239), .B(n1240), .C(n1241), .D(n1242), .S0(n1366), .S1(
        n1369), .Y(n1353) );
  MXI4XL U1209 ( .A(n1243), .B(n1244), .C(n1245), .D(n1246), .S0(n1039), .S1(
        n1373), .Y(n1304) );
  MXI4XL U1210 ( .A(n1247), .B(n1248), .C(n1249), .D(n1250), .S0(n1039), .S1(
        n1369), .Y(n1351) );
  MXI4XL U1211 ( .A(\targetX[36][3] ), .B(\targetX[38][3] ), .C(
        \targetX[37][3] ), .D(\targetX[39][3] ), .S0(n1366), .S1(n1371), .Y(
        n1349) );
  MXI4XL U1212 ( .A(\targetY[36][3] ), .B(\targetY[38][3] ), .C(
        \targetY[37][3] ), .D(\targetY[39][3] ), .S0(n1366), .S1(n1371), .Y(
        n1297) );
  MXI4XL U1213 ( .A(\targetX[32][3] ), .B(\targetX[34][3] ), .C(
        \targetX[33][3] ), .D(\targetX[35][3] ), .S0(n1366), .S1(n1371), .Y(
        n1348) );
  MXI4XL U1214 ( .A(\targetY[32][3] ), .B(\targetY[34][3] ), .C(
        \targetY[33][3] ), .D(\targetY[35][3] ), .S0(n1368), .S1(n1371), .Y(
        n1296) );
  XOR2XL U1215 ( .A(\r412/carry[5] ), .B(count[5]), .Y(N1053) );
  CLKBUFX3 U1216 ( .A(n1376), .Y(n1370) );
  OR2X4 U1217 ( .A(len1[6]), .B(len1[5]), .Y(n1390) );
  CLKBUFX3 U1218 ( .A(n1380), .Y(n1381) );
  CLKBUFX3 U1219 ( .A(n1568), .Y(n1380) );
  CLKBUFX3 U1220 ( .A(n1568), .Y(n1379) );
  CLKBUFX3 U1221 ( .A(n1568), .Y(n1378) );
  CLKINVX1 U1222 ( .A(\r401/carry[4] ), .Y(N847) );
  CLKINVX1 U1223 ( .A(\r399/carry[4] ), .Y(N830) );
  CLKBUFX3 U1224 ( .A(count[2]), .Y(n1363) );
  CLKINVX1 U1225 ( .A(N903), .Y(n1387) );
  CLKINVX1 U1226 ( .A(N903), .Y(n1383) );
  CLKBUFX3 U1227 ( .A(count[2]), .Y(n1362) );
  CLKINVX1 U1228 ( .A(\r404/carry[4] ), .Y(N952) );
  CLKINVX1 U1229 ( .A(\r406/carry[4] ), .Y(N969) );
  XNOR2X2 U1230 ( .A(n1360), .B(n1586), .Y(N965) );
  CLKINVX1 U1231 ( .A(n1065), .Y(n1385) );
  MX4X1 U1232 ( .A(\targetY[20][0] ), .B(\targetY[22][0] ), .C(
        \targetY[21][0] ), .D(\targetY[23][0] ), .S0(n1368), .S1(n1375), .Y(
        n1262) );
  MX4X1 U1233 ( .A(\targetY[4][1] ), .B(\targetY[6][1] ), .C(\targetY[5][1] ), 
        .D(\targetY[7][1] ), .S0(n1367), .S1(n1374), .Y(n1279) );
  MX4X1 U1234 ( .A(\targetY[0][1] ), .B(\targetY[2][1] ), .C(\targetY[1][1] ), 
        .D(\targetY[3][1] ), .S0(n1367), .S1(n1374), .Y(n1280) );
  MX4X1 U1235 ( .A(n1301), .B(n1299), .C(n1300), .D(n1298), .S0(n1377), .S1(
        n1363), .Y(n1302) );
  MX4X1 U1236 ( .A(\targetY[16][1] ), .B(\targetY[18][1] ), .C(
        \targetY[17][1] ), .D(\targetY[19][1] ), .S0(n1368), .S1(n1251), .Y(
        n1275) );
  MX4X1 U1237 ( .A(\targetY[24][1] ), .B(\targetY[26][1] ), .C(
        \targetY[25][1] ), .D(\targetY[27][1] ), .S0(n1368), .S1(n1251), .Y(
        n1273) );
  MX4X1 U1238 ( .A(n1288), .B(n1286), .C(n1287), .D(n1285), .S0(n1377), .S1(
        n1362), .Y(n1289) );
  MX4X1 U1239 ( .A(\targetX[12][0] ), .B(\targetX[14][0] ), .C(
        \targetX[13][0] ), .D(\targetX[15][0] ), .S0(n1367), .S1(n1373), .Y(
        n1316) );
  MX4X1 U1240 ( .A(\targetX[4][0] ), .B(\targetX[6][0] ), .C(\targetX[5][0] ), 
        .D(\targetX[7][0] ), .S0(n1367), .S1(n1373), .Y(n1318) );
  MX4X1 U1241 ( .A(\targetX[8][0] ), .B(\targetX[10][0] ), .C(\targetX[9][0] ), 
        .D(\targetX[11][0] ), .S0(n1367), .S1(n1373), .Y(n1317) );
  MX4X1 U1242 ( .A(n1358), .B(n1356), .C(n1357), .D(n1355), .S0(n1377), .S1(
        n1362), .Y(n1359) );
  MX4X1 U1243 ( .A(n1332), .B(n1330), .C(n1331), .D(n1329), .S0(n1377), .S1(
        n1363), .Y(n1333) );
  MX4X1 U1244 ( .A(n1345), .B(n1343), .C(n1344), .D(n1342), .S0(n1377), .S1(
        n1362), .Y(n1346) );
  MXI2X1 U1245 ( .A(n1296), .B(n1297), .S0(n1363), .Y(n1295) );
  MX4X1 U1246 ( .A(n1306), .B(n1304), .C(n1305), .D(n1303), .S0(n1377), .S1(
        n1363), .Y(n1307) );
  MXI2X1 U1247 ( .A(n1283), .B(n1284), .S0(n1363), .Y(n1282) );
  MX4X1 U1248 ( .A(n1293), .B(n1291), .C(n1292), .D(n1290), .S0(n1377), .S1(
        n1362), .Y(n1294) );
  MXI2X1 U1249 ( .A(n1348), .B(n1349), .S0(n1363), .Y(n1347) );
  MX4X1 U1250 ( .A(n1353), .B(n1351), .C(n1352), .D(n1350), .S0(n1377), .S1(
        n1362), .Y(n1354) );
  MXI2X1 U1251 ( .A(n1322), .B(n1323), .S0(n1363), .Y(n1321) );
  MX4X1 U1252 ( .A(n1327), .B(n1325), .C(n1326), .D(n1324), .S0(n1377), .S1(
        n1363), .Y(n1328) );
  MXI2X1 U1253 ( .A(n1335), .B(n1336), .S0(n1363), .Y(n1334) );
  MX4X1 U1254 ( .A(n1340), .B(n1338), .C(n1339), .D(n1337), .S0(n1377), .S1(
        n1362), .Y(n1341) );
  MXI4X1 U1255 ( .A(\targetY[32][1] ), .B(\targetY[34][1] ), .C(
        \targetY[33][1] ), .D(\targetY[35][1] ), .S0(n1039), .S1(n1371), .Y(
        n1270) );
  MXI4X1 U1256 ( .A(\targetY[36][1] ), .B(\targetY[38][1] ), .C(
        \targetY[37][1] ), .D(\targetY[39][1] ), .S0(n1039), .S1(n1371), .Y(
        n1271) );
  CLKINVX1 U1257 ( .A(n1098), .Y(n1388) );
  NAND2X2 U1258 ( .A(n1254), .B(n1255), .Y(\r404/carry[1] ) );
  CLKINVX1 U1259 ( .A(n1387), .Y(n1254) );
  MX4X2 U1260 ( .A(n1314), .B(n1312), .C(n1313), .D(n1311), .S0(n1377), .S1(
        n1363), .Y(n1315) );
  MXI3X2 U1261 ( .A(n1269), .B(n1264), .C(n1257), .S0(count[4]), .S1(count[5]), 
        .Y(n1360) );
  MXI3X2 U1262 ( .A(n1320), .B(n1315), .C(n1308), .S0(count[4]), .S1(count[5]), 
        .Y(n1361) );
  OAI32X2 U1263 ( .A0(n1393), .A1(len2[0]), .A2(n1392), .B0(len2[4]), .B1(
        n1392), .Y(N983) );
  OR2X8 U1264 ( .A(len2[6]), .B(len2[5]), .Y(n1392) );
  AND2X8 U1265 ( .A(n1413), .B(n1415), .Y(n1414) );
  OAI211X4 U1266 ( .A0(n1416), .A1(n1412), .B0(n1410), .C0(n1411), .Y(n1413)
         );
  XOR2X1 U1272 ( .A(\add_215/carry[5] ), .B(covered[5]), .Y(N1134) );
  OR3X1 U1273 ( .A(len1[3]), .B(len1[2]), .C(len1[1]), .Y(n1391) );
  OR3X1 U1274 ( .A(len2[3]), .B(len2[2]), .C(len2[1]), .Y(n1393) );
  OAI21XL U1275 ( .A0(n1559), .A1(n1394), .B0(n1395), .Y(n334) );
  OR3X1 U1276 ( .A(n274), .B(n1400), .C(n1401), .Y(n1399) );
  OAI21XL U1277 ( .A0(n1397), .A1(n1402), .B0(C2X[3]), .Y(n1398) );
  MXI2X1 U1278 ( .A(n1044), .B(n179), .S0(n1404), .Y(n332) );
  OAI2BB2XL U1279 ( .B0(n262), .B1(n1406), .A0N(n1382), .A1N(n1407), .Y(n331)
         );
  OAI2BB2XL U1280 ( .B0(n1047), .B1(n1406), .A0N(N1049), .A1N(n1407), .Y(n330)
         );
  OAI2BB2XL U1281 ( .B0(n260), .B1(n1406), .A0N(N1050), .A1N(n1407), .Y(n329)
         );
  OAI2BB2XL U1282 ( .B0(n259), .B1(n1406), .A0N(N1051), .A1N(n1407), .Y(n328)
         );
  OAI2BB2XL U1283 ( .B0(n258), .B1(n1406), .A0N(N1052), .A1N(n1407), .Y(n327)
         );
  OAI2BB2XL U1284 ( .B0(n257), .B1(n1406), .A0N(N1053), .A1N(n1407), .Y(n326)
         );
  AND2X1 U1285 ( .A(n1408), .B(n1409), .Y(n1407) );
  NAND3BX1 U1286 ( .AN(n1408), .B(n1410), .C(n1411), .Y(n1406) );
  OAI31XL U1287 ( .A0(n1044), .A1(state[2]), .A2(state[1]), .B0(n1412), .Y(
        n1408) );
  OAI2BB2XL U1288 ( .B0(n256), .B1(n1413), .A0N(n256), .A1N(n1414), .Y(n325)
         );
  OAI2BB2XL U1289 ( .B0(n255), .B1(n1413), .A0N(N1130), .A1N(n1414), .Y(n324)
         );
  OAI2BB2XL U1290 ( .B0(n254), .B1(n1413), .A0N(N1131), .A1N(n1414), .Y(n323)
         );
  OAI2BB2XL U1291 ( .B0(n253), .B1(n1413), .A0N(N1132), .A1N(n1414), .Y(n322)
         );
  OAI2BB2XL U1292 ( .B0(n252), .B1(n1413), .A0N(N1133), .A1N(n1414), .Y(n321)
         );
  OAI2BB2XL U1293 ( .B0(n251), .B1(n1413), .A0N(N1134), .A1N(n1414), .Y(n320)
         );
  NAND3BX1 U1294 ( .AN(n248), .B(n1421), .C(n1422), .Y(n1420) );
  OAI21XL U1295 ( .A0(n1422), .A1(n1423), .B0(C2Y[3]), .Y(n1419) );
  OAI21XL U1296 ( .A0(n1558), .A1(n1394), .B0(n1425), .Y(n316) );
  MXI2X1 U1297 ( .A(n1402), .B(n1426), .S0(n275), .Y(n1425) );
  NOR2X1 U1298 ( .A(n276), .B(n1401), .Y(n1426) );
  OAI21XL U1299 ( .A0(n1557), .A1(n1394), .B0(n1427), .Y(n314) );
  MXI2X1 U1300 ( .A(n1428), .B(n1429), .S0(n274), .Y(n1427) );
  NOR2X1 U1301 ( .A(n1400), .B(n1401), .Y(n1429) );
  CLKINVX1 U1302 ( .A(n1432), .Y(n1396) );
  NAND2X1 U1303 ( .A(n1434), .B(n1435), .Y(n1432) );
  OAI21XL U1304 ( .A0(n1405), .A1(n1436), .B0(n1437), .Y(n1435) );
  OAI21XL U1305 ( .A0(n1554), .A1(n1418), .B0(n1438), .Y(n313) );
  OAI21XL U1306 ( .A0(n1418), .A1(n1441), .B0(n1442), .Y(n311) );
  MXI2X1 U1307 ( .A(n1443), .B(n1444), .S0(n249), .Y(n1442) );
  NOR2X1 U1308 ( .A(n250), .B(n1440), .Y(n1444) );
  OAI21XL U1309 ( .A0(n1553), .A1(n1418), .B0(n1445), .Y(n309) );
  MXI2X1 U1310 ( .A(n1423), .B(n1446), .S0(n248), .Y(n1445) );
  NOR2X1 U1311 ( .A(n1447), .B(n1440), .Y(n1446) );
  CLKINVX1 U1312 ( .A(n1422), .Y(n1440) );
  AO21X1 U1313 ( .A0(n1422), .A1(n249), .B0(n1443), .Y(n1423) );
  NOR2X1 U1314 ( .A(n1431), .B(n1436), .Y(n1422) );
  CLKINVX1 U1315 ( .A(n1449), .Y(n1448) );
  OAI21XL U1316 ( .A0(n251), .A1(n1450), .B0(n187), .Y(n302) );
  NAND2X1 U1317 ( .A(n1451), .B(n1449), .Y(n301) );
  NOR2X1 U1318 ( .A(n1454), .B(n1455), .Y(n1453) );
  OAI221XL U1319 ( .A0(n271), .A1(n1457), .B0(n1560), .B1(n1458), .C0(n1459), 
        .Y(n299) );
  OAI21XL U1320 ( .A0(n1460), .A1(n1461), .B0(C1Y[3]), .Y(n1459) );
  CLKINVX1 U1321 ( .A(n1463), .Y(n1457) );
  OAI21XL U1322 ( .A0(n1468), .A1(n1469), .B0(C1X[3]), .Y(n1465) );
  OAI21XL U1323 ( .A0(n1563), .A1(n1464), .B0(n1471), .Y(n296) );
  OAI21XL U1324 ( .A0(n1562), .A1(n1464), .B0(n1473), .Y(n294) );
  MXI2X1 U1325 ( .A(n1469), .B(n1474), .S0(n268), .Y(n1473) );
  NOR2X1 U1326 ( .A(n269), .B(n1475), .Y(n1474) );
  OAI21XL U1327 ( .A0(n1561), .A1(n1464), .B0(n1476), .Y(n292) );
  MXI2X1 U1328 ( .A(n1477), .B(n1478), .S0(n267), .Y(n1476) );
  NOR2X1 U1329 ( .A(n1479), .B(n1475), .Y(n1478) );
  CLKINVX1 U1330 ( .A(n1480), .Y(n1472) );
  OAI2BB1X1 U1331 ( .A0N(n1433), .A1N(n1482), .B0(n1483), .Y(n1480) );
  OAI21XL U1332 ( .A0(n1566), .A1(n1458), .B0(n1484), .Y(n291) );
  CLKMX2X2 U1333 ( .A(n1485), .B(n1486), .S0(n273), .Y(n1484) );
  OAI21XL U1334 ( .A0(n1458), .A1(n1487), .B0(n1488), .Y(n289) );
  MXI2X1 U1335 ( .A(n1461), .B(n1489), .S0(n272), .Y(n1488) );
  NOR2X1 U1336 ( .A(n273), .B(n1486), .Y(n1489) );
  OAI21XL U1337 ( .A0(n1565), .A1(n1458), .B0(n1490), .Y(n287) );
  MXI2X1 U1338 ( .A(n1491), .B(n1463), .S0(n271), .Y(n1490) );
  NOR3X1 U1339 ( .A(n272), .B(n273), .C(n1486), .Y(n1463) );
  CLKINVX1 U1340 ( .A(n1460), .Y(n1486) );
  AO21X1 U1341 ( .A0(n1460), .A1(n272), .B0(n1461), .Y(n1491) );
  OAI2BB1X1 U1342 ( .A0N(n1460), .A1N(n273), .B0(n1485), .Y(n1461) );
  NOR2X1 U1343 ( .A(n1410), .B(n1482), .Y(n1460) );
  NOR2X1 U1344 ( .A(n1493), .B(state[0]), .Y(n1433) );
  CLKINVX1 U1345 ( .A(n1454), .Y(n1431) );
  CLKINVX1 U1346 ( .A(n1411), .Y(n1437) );
  NOR2X1 U1347 ( .A(n1405), .B(n1454), .Y(n1411) );
  OAI21XL U1348 ( .A0(n251), .A1(n1496), .B0(n202), .Y(n278) );
  OAI221XL U1349 ( .A0(n1498), .A1(n1499), .B0(n251), .B1(n1500), .C0(n1501), 
        .Y(n1497) );
  NAND3X1 U1350 ( .A(n1502), .B(covered[4]), .C(n201), .Y(n1501) );
  OAI21XL U1351 ( .A0(n201), .A1(covered[4]), .B0(n1502), .Y(n1499) );
  NAND2X1 U1352 ( .A(n251), .B(n1500), .Y(n1502) );
  AOI22X1 U1353 ( .A0(n1503), .A1(covered[3]), .B0(n1504), .B1(n200), .Y(n1498) );
  OR2X1 U1354 ( .A(n1504), .B(n200), .Y(n1503) );
  OAI2BB1X1 U1355 ( .A0N(n1505), .A1N(n199), .B0(n1506), .Y(n1504) );
  OAI21XL U1356 ( .A0(n199), .A1(n1505), .B0(covered[2]), .Y(n1506) );
  OAI2BB1X1 U1357 ( .A0N(covered[1]), .A1N(n198), .B0(n1507), .Y(n1505) );
  OAI22XL U1358 ( .A0(n197), .A1(covered[0]), .B0(n198), .B1(covered[1]), .Y(
        n1507) );
  OAI221XL U1359 ( .A0(n1510), .A1(n1511), .B0(n251), .B1(n1512), .C0(n1513), 
        .Y(n1508) );
  NAND3X1 U1360 ( .A(n1514), .B(covered[4]), .C(n186), .Y(n1513) );
  OAI21XL U1361 ( .A0(n186), .A1(covered[4]), .B0(n1514), .Y(n1511) );
  NAND2X1 U1362 ( .A(n251), .B(n1512), .Y(n1514) );
  AOI2BB2X1 U1363 ( .B0(n1515), .B1(covered[3]), .A0N(n1516), .A1N(n1517), .Y(
        n1510) );
  NAND2X1 U1364 ( .A(n1516), .B(n1517), .Y(n1515) );
  ACHCONX2 U1365 ( .A(covered[2]), .B(n1518), .CI(n263), .CON(n1517) );
  OAI2BB1X1 U1366 ( .A0N(covered[1]), .A1N(n264), .B0(n1519), .Y(n1518) );
  OAI22XL U1367 ( .A0(n265), .A1(covered[0]), .B0(n264), .B1(covered[1]), .Y(
        n1519) );
  NAND2X1 U1368 ( .A(n1509), .B(n1449), .Y(n245) );
  NAND3X1 U1369 ( .A(n1454), .B(n1436), .C(n1430), .Y(n1449) );
  NOR3X1 U1370 ( .A(n204), .B(n274), .C(n1400), .Y(n1430) );
  OR2X1 U1371 ( .A(n275), .B(n276), .Y(n1400) );
  NOR2X1 U1372 ( .A(n1044), .B(n1493), .Y(n1454) );
  NAND3X1 U1373 ( .A(n1366), .B(n1374), .C(n260), .Y(n1527) );
  NAND3X1 U1374 ( .A(n1362), .B(n1374), .C(n1047), .Y(n1529) );
  NAND3X1 U1375 ( .A(n260), .B(n1374), .C(n1047), .Y(n1530) );
  NAND3X1 U1376 ( .A(n1362), .B(n1367), .C(n262), .Y(n1531) );
  NAND3X1 U1377 ( .A(n1047), .B(n1362), .C(n262), .Y(n1532) );
  NAND3X1 U1378 ( .A(n260), .B(n1367), .C(n262), .Y(n1533) );
  NAND3X1 U1379 ( .A(n1047), .B(n260), .C(n262), .Y(n1534) );
  AND2X1 U1380 ( .A(n257), .B(n1520), .Y(n1535) );
  NOR4X1 U1381 ( .A(n1044), .B(RST), .C(state[1]), .D(state[2]), .Y(n1520) );
  OAI211X1 U1382 ( .A0(n1536), .A1(n1412), .B0(n1537), .C0(n1493), .Y(N1023)
         );
  NAND2X1 U1383 ( .A(state[1]), .B(n1045), .Y(n1493) );
  CLKINVX1 U1384 ( .A(n1538), .Y(n1536) );
  NOR2X1 U1385 ( .A(n1412), .B(n1538), .Y(N1022) );
  OAI31XL U1386 ( .A0(n1521), .A1(state[2]), .A2(state[1]), .B0(n1541), .Y(
        N1021) );
  NAND4X1 U1387 ( .A(n185), .B(n263), .C(n265), .D(n1543), .Y(n1539) );
  AND3X1 U1388 ( .A(n264), .B(n187), .C(n186), .Y(n1543) );
  OAI21XL U1389 ( .A0(n1409), .A1(n1544), .B0(n1540), .Y(n1542) );
  NAND4X1 U1390 ( .A(n1545), .B(n1546), .C(n1547), .D(n1548), .Y(n1540) );
  NOR3X1 U1391 ( .A(n1549), .B(n1550), .C(n1551), .Y(n1548) );
  XNOR2X1 U1392 ( .A(n200), .B(n1516), .Y(n1551) );
  XNOR2X1 U1393 ( .A(n1500), .B(n187), .Y(n1550) );
  XOR2X1 U1394 ( .A(n201), .B(n186), .Y(n1549) );
  XNOR2X1 U1395 ( .A(n198), .B(n264), .Y(n1547) );
  XNOR2X1 U1396 ( .A(n199), .B(n263), .Y(n1546) );
  XNOR2X1 U1397 ( .A(n197), .B(n265), .Y(n1545) );
  MXI2X1 U1398 ( .A(n1492), .B(n1434), .S0(n1455), .Y(n1544) );
  NAND4X1 U1399 ( .A(n276), .B(n275), .C(n1552), .D(n274), .Y(n1434) );
  NOR2BX1 U1400 ( .AN(n1436), .B(C2X[3]), .Y(n1552) );
  NOR3X1 U1401 ( .A(n247), .B(n248), .C(n1447), .Y(n1436) );
  CLKINVX1 U1402 ( .A(n1421), .Y(n1447) );
  NOR2X1 U1403 ( .A(n249), .B(n250), .Y(n1421) );
  CLKINVX1 U1404 ( .A(n1452), .Y(n1492) );
  NAND2X1 U1405 ( .A(n1481), .B(n1482), .Y(n1452) );
  NOR4X1 U1406 ( .A(n270), .B(n271), .C(n272), .D(n273), .Y(n1482) );
  NOR3X1 U1407 ( .A(n266), .B(n267), .C(n1479), .Y(n1481) );
  CLKINVX1 U1408 ( .A(n1467), .Y(n1479) );
  NOR2X1 U1409 ( .A(n268), .B(n269), .Y(n1467) );
  NAND3X1 U1410 ( .A(n1366), .B(n1374), .C(n1362), .Y(n1522) );
  NAND2X1 U1411 ( .A(state[2]), .B(state[1]), .Y(N1020) );
endmodule

